// Verilog pattern output written by  TetraMAX (TM)  B-2008.09-SP2-i081128_181834 
// Date: Wed Jul  6 12:09:50 2011
// Module tested: c7552

//     Uncollapsed Stuck Fault Summary Report
// -----------------------------------------------
// fault class                     code   #faults
// ------------------------------  ----  ---------
// Detected                         DT       6578
// Possibly detected                PT          0
// Undetectable                     UD          0
// ATPG untestable                  AU          0
// Not detected                     ND        310
// -----------------------------------------------
// total faults                              6888
// test coverage                            95.50%
// -----------------------------------------------
// 
//            Pattern Summary Report
// -----------------------------------------------
// #internal patterns                         181
//     #basic_scan patterns                   181
// -----------------------------------------------
// 
// There are no rule fails
// There are no clocks
// There are no constraint ports
// There are no equivalent pins
// There are no net connections

`timescale 1 ns / 1 ns

//
// --- NOTE: Remove the comment to define 'tmax_iddq' to activate processing of IDDQ events
//     Or use '+define+tmax_iddq' on the verilog compile line
//
//`define tmax_iddq

module AAA_tmax_testbench_1_16 ;
   parameter NAMELENGTH = 200; // max length of names reported in fails
   integer nofails, bit, pattern, lastpattern;
   integer error_banner; // flag for tracking displayed error banner
   integer loads;        // number of load_unloads for current pattern
   integer patm1;        // pattern - 1
   integer patp1;        // pattern + lastpattern
   integer prev_pat;     // previous pattern number
   integer report_interval; // report pattern progress every Nth pattern
   integer verbose;      // message verbosity level
   parameter NINPUTS = 207, NOUTPUTS = 108;
   wire [0:NOUTPUTS-1] PO; reg [0:NOUTPUTS-1] ALLPOS, XPCT, MASK;
   reg [0:NINPUTS-1] PI, ALLPIS;
   reg [0:8*(NAMELENGTH-1)] POnames [0:NOUTPUTS-1];
   event IDDQ;

   wire N1;
   wire N5;
   wire N9;
   wire N12;
   wire N15;
   wire N18;
   wire N23;
   wire N26;
   wire N29;
   wire N32;
   wire N35;
   wire N38;
   wire N41;
   wire N44;
   wire N47;
   wire N50;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N69;
   wire N70;
   wire N73;
   wire N74;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N82;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N94;
   wire N97;
   wire N100;
   wire N103;
   wire N106;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N118;
   wire N121;
   wire N124;
   wire N127;
   wire N130;
   wire N133;
   wire N134;
   wire N135;
   wire N138;
   wire N141;
   wire N144;
   wire N147;
   wire N150;
   wire N151;
   wire N152;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N178;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire N185;
   wire N186;
   wire N187;
   wire N188;
   wire N189;
   wire N190;
   wire N191;
   wire N192;
   wire N193;
   wire N194;
   wire N195;
   wire N196;
   wire N197;
   wire N198;
   wire N199;
   wire N200;
   wire N201;
   wire N202;
   wire N203;
   wire N204;
   wire N205;
   wire N206;
   wire N207;
   wire N208;
   wire N209;
   wire N210;
   wire N211;
   wire N212;
   wire N213;
   wire N214;
   wire N215;
   wire N216;
   wire N217;
   wire N218;
   wire N219;
   wire N220;
   wire N221;
   wire N222;
   wire N223;
   wire N224;
   wire N225;
   wire N226;
   wire N227;
   wire N228;
   wire N229;
   wire N230;
   wire N231;
   wire N232;
   wire N233;
   wire N234;
   wire N235;
   wire N236;
   wire N237;
   wire N238;
   wire N239;
   wire N240;
   wire N242;
   wire N245;
   wire N248;
   wire N251;
   wire N254;
   wire N257;
   wire N260;
   wire N263;
   wire N267;
   wire N271;
   wire N274;
   wire N277;
   wire N280;
   wire N283;
   wire N286;
   wire N289;
   wire N293;
   wire N296;
   wire N299;
   wire N303;
   wire N307;
   wire N310;
   wire N313;
   wire N316;
   wire N319;
   wire N322;
   wire N325;
   wire N328;
   wire N331;
   wire N334;
   wire N337;
   wire N340;
   wire N343;
   wire N346;
   wire N349;
   wire N352;
   wire N355;
   wire N358;
   wire N361;
   wire N364;
   wire N367;
   wire N382;
   wire N241_I;
   wire N387;
   wire N388;
   wire N478;
   wire N482;
   wire N484;
   wire N486;
   wire N489;
   wire N492;
   wire N501;
   wire N505;
   wire N507;
   wire N509;
   wire N511;
   wire N513;
   wire N515;
   wire N517;
   wire N519;
   wire N535;
   wire N537;
   wire N539;
   wire N541;
   wire N543;
   wire N545;
   wire N547;
   wire N549;
   wire N551;
   wire N553;
   wire N556;
   wire N559;
   wire N561;
   wire N563;
   wire N565;
   wire N567;
   wire N569;
   wire N571;
   wire N573;
   wire N582;
   wire N643;
   wire N707;
   wire N813;
   wire N881;
   wire N882;
   wire N883;
   wire N884;
   wire N885;
   wire N889;
   wire N945;
   wire N1110;
   wire N1111;
   wire N1112;
   wire N1113;
   wire N1114;
   wire N1489;
   wire N1490;
   wire N1781;
   wire N10025;
   wire N10101;
   wire N10102;
   wire N10103;
   wire N10104;
   wire N10109;
   wire N10110;
   wire N10111;
   wire N10112;
   wire N10350;
   wire N10351;
   wire N10352;
   wire N10353;
   wire N10574;
   wire N10575;
   wire N10576;
   wire N10628;
   wire N10632;
   wire N10641;
   wire N10704;
   wire N10706;
   wire N10711;
   wire N10712;
   wire N10713;
   wire N10714;
   wire N10715;
   wire N10716;
   wire N10717;
   wire N10718;
   wire N10729;
   wire N10759;
   wire N10760;
   wire N10761;
   wire N10762;
   wire N10763;
   wire N10827;
   wire N10837;
   wire N10838;
   wire N10839;
   wire N10840;
   wire N10868;
   wire N10869;
   wire N10870;
   wire N10871;
   wire N10905;
   wire N10906;
   wire N10907;
   wire N10908;
   wire N11333;
   wire N11334;
   wire N11340;
   wire N11342;
   wire N241_O;

   // map PI[] vector to DUT inputs and bidis
   assign N1 = PI[0];
   assign N5 = PI[1];
   assign N9 = PI[2];
   assign N12 = PI[3];
   assign N15 = PI[4];
   assign N18 = PI[5];
   assign N23 = PI[6];
   assign N26 = PI[7];
   assign N29 = PI[8];
   assign N32 = PI[9];
   assign N35 = PI[10];
   assign N38 = PI[11];
   assign N41 = PI[12];
   assign N44 = PI[13];
   assign N47 = PI[14];
   assign N50 = PI[15];
   assign N53 = PI[16];
   assign N54 = PI[17];
   assign N55 = PI[18];
   assign N56 = PI[19];
   assign N57 = PI[20];
   assign N58 = PI[21];
   assign N59 = PI[22];
   assign N60 = PI[23];
   assign N61 = PI[24];
   assign N62 = PI[25];
   assign N63 = PI[26];
   assign N64 = PI[27];
   assign N65 = PI[28];
   assign N66 = PI[29];
   assign N69 = PI[30];
   assign N70 = PI[31];
   assign N73 = PI[32];
   assign N74 = PI[33];
   assign N75 = PI[34];
   assign N76 = PI[35];
   assign N77 = PI[36];
   assign N78 = PI[37];
   assign N79 = PI[38];
   assign N80 = PI[39];
   assign N81 = PI[40];
   assign N82 = PI[41];
   assign N83 = PI[42];
   assign N84 = PI[43];
   assign N85 = PI[44];
   assign N86 = PI[45];
   assign N87 = PI[46];
   assign N88 = PI[47];
   assign N89 = PI[48];
   assign N94 = PI[49];
   assign N97 = PI[50];
   assign N100 = PI[51];
   assign N103 = PI[52];
   assign N106 = PI[53];
   assign N109 = PI[54];
   assign N110 = PI[55];
   assign N111 = PI[56];
   assign N112 = PI[57];
   assign N113 = PI[58];
   assign N114 = PI[59];
   assign N115 = PI[60];
   assign N118 = PI[61];
   assign N121 = PI[62];
   assign N124 = PI[63];
   assign N127 = PI[64];
   assign N130 = PI[65];
   assign N133 = PI[66];
   assign N134 = PI[67];
   assign N135 = PI[68];
   assign N138 = PI[69];
   assign N141 = PI[70];
   assign N144 = PI[71];
   assign N147 = PI[72];
   assign N150 = PI[73];
   assign N151 = PI[74];
   assign N152 = PI[75];
   assign N153 = PI[76];
   assign N154 = PI[77];
   assign N155 = PI[78];
   assign N156 = PI[79];
   assign N157 = PI[80];
   assign N158 = PI[81];
   assign N159 = PI[82];
   assign N160 = PI[83];
   assign N161 = PI[84];
   assign N162 = PI[85];
   assign N163 = PI[86];
   assign N164 = PI[87];
   assign N165 = PI[88];
   assign N166 = PI[89];
   assign N167 = PI[90];
   assign N168 = PI[91];
   assign N169 = PI[92];
   assign N170 = PI[93];
   assign N171 = PI[94];
   assign N172 = PI[95];
   assign N173 = PI[96];
   assign N174 = PI[97];
   assign N175 = PI[98];
   assign N176 = PI[99];
   assign N177 = PI[100];
   assign N178 = PI[101];
   assign N179 = PI[102];
   assign N180 = PI[103];
   assign N181 = PI[104];
   assign N182 = PI[105];
   assign N183 = PI[106];
   assign N184 = PI[107];
   assign N185 = PI[108];
   assign N186 = PI[109];
   assign N187 = PI[110];
   assign N188 = PI[111];
   assign N189 = PI[112];
   assign N190 = PI[113];
   assign N191 = PI[114];
   assign N192 = PI[115];
   assign N193 = PI[116];
   assign N194 = PI[117];
   assign N195 = PI[118];
   assign N196 = PI[119];
   assign N197 = PI[120];
   assign N198 = PI[121];
   assign N199 = PI[122];
   assign N200 = PI[123];
   assign N201 = PI[124];
   assign N202 = PI[125];
   assign N203 = PI[126];
   assign N204 = PI[127];
   assign N205 = PI[128];
   assign N206 = PI[129];
   assign N207 = PI[130];
   assign N208 = PI[131];
   assign N209 = PI[132];
   assign N210 = PI[133];
   assign N211 = PI[134];
   assign N212 = PI[135];
   assign N213 = PI[136];
   assign N214 = PI[137];
   assign N215 = PI[138];
   assign N216 = PI[139];
   assign N217 = PI[140];
   assign N218 = PI[141];
   assign N219 = PI[142];
   assign N220 = PI[143];
   assign N221 = PI[144];
   assign N222 = PI[145];
   assign N223 = PI[146];
   assign N224 = PI[147];
   assign N225 = PI[148];
   assign N226 = PI[149];
   assign N227 = PI[150];
   assign N228 = PI[151];
   assign N229 = PI[152];
   assign N230 = PI[153];
   assign N231 = PI[154];
   assign N232 = PI[155];
   assign N233 = PI[156];
   assign N234 = PI[157];
   assign N235 = PI[158];
   assign N236 = PI[159];
   assign N237 = PI[160];
   assign N238 = PI[161];
   assign N239 = PI[162];
   assign N240 = PI[163];
   assign N242 = PI[164];
   assign N245 = PI[165];
   assign N248 = PI[166];
   assign N251 = PI[167];
   assign N254 = PI[168];
   assign N257 = PI[169];
   assign N260 = PI[170];
   assign N263 = PI[171];
   assign N267 = PI[172];
   assign N271 = PI[173];
   assign N274 = PI[174];
   assign N277 = PI[175];
   assign N280 = PI[176];
   assign N283 = PI[177];
   assign N286 = PI[178];
   assign N289 = PI[179];
   assign N293 = PI[180];
   assign N296 = PI[181];
   assign N299 = PI[182];
   assign N303 = PI[183];
   assign N307 = PI[184];
   assign N310 = PI[185];
   assign N313 = PI[186];
   assign N316 = PI[187];
   assign N319 = PI[188];
   assign N322 = PI[189];
   assign N325 = PI[190];
   assign N328 = PI[191];
   assign N331 = PI[192];
   assign N334 = PI[193];
   assign N337 = PI[194];
   assign N340 = PI[195];
   assign N343 = PI[196];
   assign N346 = PI[197];
   assign N349 = PI[198];
   assign N352 = PI[199];
   assign N355 = PI[200];
   assign N358 = PI[201];
   assign N361 = PI[202];
   assign N364 = PI[203];
   assign N367 = PI[204];
   assign N382 = PI[205];
   assign N241_I = PI[206];

   // map DUT outputs and bidis to PO[] vector
   assign
      PO[0] = N387 ,
      PO[1] = N388 ,
      PO[2] = N478 ,
      PO[3] = N482 ,
      PO[4] = N484 ,
      PO[5] = N486 ,
      PO[6] = N489 ,
      PO[7] = N492 ,
      PO[8] = N501 ,
      PO[9] = N505 ,
      PO[10] = N507 ,
      PO[11] = N509 ,
      PO[12] = N511 ,
      PO[13] = N513 ,
      PO[14] = N515 ,
      PO[15] = N517 ,
      PO[16] = N519 ,
      PO[17] = N535 ,
      PO[18] = N537 ,
      PO[19] = N539 ,
      PO[20] = N541 ,
      PO[21] = N543 ,
      PO[22] = N545 ,
      PO[23] = N547 ,
      PO[24] = N549 ,
      PO[25] = N551 ,
      PO[26] = N553 ,
      PO[27] = N556 ,
      PO[28] = N559 ,
      PO[29] = N561 ,
      PO[30] = N563 ,
      PO[31] = N565 ;
   assign
      PO[32] = N567 ,
      PO[33] = N569 ,
      PO[34] = N571 ,
      PO[35] = N573 ,
      PO[36] = N582 ,
      PO[37] = N643 ,
      PO[38] = N707 ,
      PO[39] = N813 ,
      PO[40] = N881 ,
      PO[41] = N882 ,
      PO[42] = N883 ,
      PO[43] = N884 ,
      PO[44] = N885 ,
      PO[45] = N889 ,
      PO[46] = N945 ,
      PO[47] = N1110 ,
      PO[48] = N1111 ,
      PO[49] = N1112 ,
      PO[50] = N1113 ,
      PO[51] = N1114 ,
      PO[52] = N1489 ,
      PO[53] = N1490 ,
      PO[54] = N1781 ,
      PO[55] = N10025 ,
      PO[56] = N10101 ,
      PO[57] = N10102 ,
      PO[58] = N10103 ,
      PO[59] = N10104 ,
      PO[60] = N10109 ,
      PO[61] = N10110 ,
      PO[62] = N10111 ,
      PO[63] = N10112 ;
   assign
      PO[64] = N10350 ,
      PO[65] = N10351 ,
      PO[66] = N10352 ,
      PO[67] = N10353 ,
      PO[68] = N10574 ,
      PO[69] = N10575 ,
      PO[70] = N10576 ,
      PO[71] = N10628 ,
      PO[72] = N10632 ,
      PO[73] = N10641 ,
      PO[74] = N10704 ,
      PO[75] = N10706 ,
      PO[76] = N10711 ,
      PO[77] = N10712 ,
      PO[78] = N10713 ,
      PO[79] = N10714 ,
      PO[80] = N10715 ,
      PO[81] = N10716 ,
      PO[82] = N10717 ,
      PO[83] = N10718 ,
      PO[84] = N10729 ,
      PO[85] = N10759 ,
      PO[86] = N10760 ,
      PO[87] = N10761 ,
      PO[88] = N10762 ,
      PO[89] = N10763 ,
      PO[90] = N10827 ,
      PO[91] = N10837 ,
      PO[92] = N10838 ,
      PO[93] = N10839 ,
      PO[94] = N10840 ,
      PO[95] = N10868 ;
   assign
      PO[96] = N10869 ,
      PO[97] = N10870 ,
      PO[98] = N10871 ,
      PO[99] = N10905 ,
      PO[100] = N10906 ,
      PO[101] = N10907 ,
      PO[102] = N10908 ,
      PO[103] = N11333 ,
      PO[104] = N11334 ,
      PO[105] = N11340 ,
      PO[106] = N11342 ,
      PO[107] = N241_O ;

   // instantiate the design into the testbench
   c7552 dut (
      .N1(N1),
      .N5(N5),
      .N9(N9),
      .N12(N12),
      .N15(N15),
      .N18(N18),
      .N23(N23),
      .N26(N26),
      .N29(N29),
      .N32(N32),
      .N35(N35),
      .N38(N38),
      .N41(N41),
      .N44(N44),
      .N47(N47),
      .N50(N50),
      .N53(N53),
      .N54(N54),
      .N55(N55),
      .N56(N56),
      .N57(N57),
      .N58(N58),
      .N59(N59),
      .N60(N60),
      .N61(N61),
      .N62(N62),
      .N63(N63),
      .N64(N64),
      .N65(N65),
      .N66(N66),
      .N69(N69),
      .N70(N70),
      .N73(N73),
      .N74(N74),
      .N75(N75),
      .N76(N76),
      .N77(N77),
      .N78(N78),
      .N79(N79),
      .N80(N80),
      .N81(N81),
      .N82(N82),
      .N83(N83),
      .N84(N84),
      .N85(N85),
      .N86(N86),
      .N87(N87),
      .N88(N88),
      .N89(N89),
      .N94(N94),
      .N97(N97),
      .N100(N100),
      .N103(N103),
      .N106(N106),
      .N109(N109),
      .N110(N110),
      .N111(N111),
      .N112(N112),
      .N113(N113),
      .N114(N114),
      .N115(N115),
      .N118(N118),
      .N121(N121),
      .N124(N124),
      .N127(N127),
      .N130(N130),
      .N133(N133),
      .N134(N134),
      .N135(N135),
      .N138(N138),
      .N141(N141),
      .N144(N144),
      .N147(N147),
      .N150(N150),
      .N151(N151),
      .N152(N152),
      .N153(N153),
      .N154(N154),
      .N155(N155),
      .N156(N156),
      .N157(N157),
      .N158(N158),
      .N159(N159),
      .N160(N160),
      .N161(N161),
      .N162(N162),
      .N163(N163),
      .N164(N164),
      .N165(N165),
      .N166(N166),
      .N167(N167),
      .N168(N168),
      .N169(N169),
      .N170(N170),
      .N171(N171),
      .N172(N172),
      .N173(N173),
      .N174(N174),
      .N175(N175),
      .N176(N176),
      .N177(N177),
      .N178(N178),
      .N179(N179),
      .N180(N180),
      .N181(N181),
      .N182(N182),
      .N183(N183),
      .N184(N184),
      .N185(N185),
      .N186(N186),
      .N187(N187),
      .N188(N188),
      .N189(N189),
      .N190(N190),
      .N191(N191),
      .N192(N192),
      .N193(N193),
      .N194(N194),
      .N195(N195),
      .N196(N196),
      .N197(N197),
      .N198(N198),
      .N199(N199),
      .N200(N200),
      .N201(N201),
      .N202(N202),
      .N203(N203),
      .N204(N204),
      .N205(N205),
      .N206(N206),
      .N207(N207),
      .N208(N208),
      .N209(N209),
      .N210(N210),
      .N211(N211),
      .N212(N212),
      .N213(N213),
      .N214(N214),
      .N215(N215),
      .N216(N216),
      .N217(N217),
      .N218(N218),
      .N219(N219),
      .N220(N220),
      .N221(N221),
      .N222(N222),
      .N223(N223),
      .N224(N224),
      .N225(N225),
      .N226(N226),
      .N227(N227),
      .N228(N228),
      .N229(N229),
      .N230(N230),
      .N231(N231),
      .N232(N232),
      .N233(N233),
      .N234(N234),
      .N235(N235),
      .N236(N236),
      .N237(N237),
      .N238(N238),
      .N239(N239),
      .N240(N240),
      .N242(N242),
      .N245(N245),
      .N248(N248),
      .N251(N251),
      .N254(N254),
      .N257(N257),
      .N260(N260),
      .N263(N263),
      .N267(N267),
      .N271(N271),
      .N274(N274),
      .N277(N277),
      .N280(N280),
      .N283(N283),
      .N286(N286),
      .N289(N289),
      .N293(N293),
      .N296(N296),
      .N299(N299),
      .N303(N303),
      .N307(N307),
      .N310(N310),
      .N313(N313),
      .N316(N316),
      .N319(N319),
      .N322(N322),
      .N325(N325),
      .N328(N328),
      .N331(N331),
      .N334(N334),
      .N337(N337),
      .N340(N340),
      .N343(N343),
      .N346(N346),
      .N349(N349),
      .N352(N352),
      .N355(N355),
      .N358(N358),
      .N361(N361),
      .N364(N364),
      .N367(N367),
      .N382(N382),
      .N241_I(N241_I),
      .N387(N387),
      .N388(N388),
      .N478(N478),
      .N482(N482),
      .N484(N484),
      .N486(N486),
      .N489(N489),
      .N492(N492),
      .N501(N501),
      .N505(N505),
      .N507(N507),
      .N509(N509),
      .N511(N511),
      .N513(N513),
      .N515(N515),
      .N517(N517),
      .N519(N519),
      .N535(N535),
      .N537(N537),
      .N539(N539),
      .N541(N541),
      .N543(N543),
      .N545(N545),
      .N547(N547),
      .N549(N549),
      .N551(N551),
      .N553(N553),
      .N556(N556),
      .N559(N559),
      .N561(N561),
      .N563(N563),
      .N565(N565),
      .N567(N567),
      .N569(N569),
      .N571(N571),
      .N573(N573),
      .N582(N582),
      .N643(N643),
      .N707(N707),
      .N813(N813),
      .N881(N881),
      .N882(N882),
      .N883(N883),
      .N884(N884),
      .N885(N885),
      .N889(N889),
      .N945(N945),
      .N1110(N1110),
      .N1111(N1111),
      .N1112(N1112),
      .N1113(N1113),
      .N1114(N1114),
      .N1489(N1489),
      .N1490(N1490),
      .N1781(N1781),
      .N10025(N10025),
      .N10101(N10101),
      .N10102(N10102),
      .N10103(N10103),
      .N10104(N10104),
      .N10109(N10109),
      .N10110(N10110),
      .N10111(N10111),
      .N10112(N10112),
      .N10350(N10350),
      .N10351(N10351),
      .N10352(N10352),
      .N10353(N10353),
      .N10574(N10574),
      .N10575(N10575),
      .N10576(N10576),
      .N10628(N10628),
      .N10632(N10632),
      .N10641(N10641),
      .N10704(N10704),
      .N10706(N10706),
      .N10711(N10711),
      .N10712(N10712),
      .N10713(N10713),
      .N10714(N10714),
      .N10715(N10715),
      .N10716(N10716),
      .N10717(N10717),
      .N10718(N10718),
      .N10729(N10729),
      .N10759(N10759),
      .N10760(N10760),
      .N10761(N10761),
      .N10762(N10762),
      .N10763(N10763),
      .N10827(N10827),
      .N10837(N10837),
      .N10838(N10838),
      .N10839(N10839),
      .N10840(N10840),
      .N10868(N10868),
      .N10869(N10869),
      .N10870(N10870),
      .N10871(N10871),
      .N10905(N10905),
      .N10906(N10906),
      .N10907(N10907),
      .N10908(N10908),
      .N11333(N11333),
      .N11334(N11334),
      .N11340(N11340),
      .N11342(N11342),
      .N241_O(N241_O)   );


   integer errshown;
   event measurePO;
   always @ measurePO begin
      if (((XPCT&MASK) !== (ALLPOS&MASK)) || (XPCT !== (~(~XPCT)))) begin
         errshown = 0;
         for (bit = 0; bit < NOUTPUTS; bit=bit + 1) begin
            if (MASK[bit]==1'b1) begin
               if (XPCT[bit] !== ALLPOS[bit]) begin
                  if (errshown==0) $display("\n// *** ERROR during capture pattern %0d, T=%t", pattern, $time);
                  $display("  %0d %0s (exp=%b, got=%b)", pattern, POnames[bit], XPCT[bit], ALLPOS[bit]);
                  nofails = nofails + 1; errshown = 1;
               end
            end
         end
      end
   end

   event forcePI_default_WFT;
   always @ forcePI_default_WFT begin
      PI = ALLPIS;
   end
   event measurePO_default_WFT;
   always @ measurePO_default_WFT begin
      #40;
      ALLPOS = PO;
      #0; #0 -> measurePO;
      `ifdef tmax_iddq
         #0; ->IDDQ;
      `endif
   end

   always @ IDDQ begin
   `ifdef tmax_iddq
      $ssi_iddq("strobe_try");
      $ssi_iddq("status drivers leaky AAA_tmax_testbench_1_16.leaky");
   `endif
   end

   event capture;
   always @ capture begin
      ->forcePI_default_WFT;
      #100; ->measurePO_default_WFT;
   end


   initial begin

      //
      // --- establish a default time format for %t
      //
      $timeformat(-9,2," ns",18);

      //
      // --- default verbosity to 2 but also allow user override by
      //     using '+define+tmax_msg=N' on verilog compile line.
      //
      `ifdef tmax_msg
         verbose = `tmax_msg ;
      `else
         verbose = 2 ;
      `endif

      //
      // --- default pattern reporting interval to 5 but also allow user
      //     override by using '+define+tmax_rpt=N' on verilog compile line.
      //
      `ifdef tmax_rpt
         report_interval = `tmax_rpt ;
      `else
         report_interval = 5 ;
      `endif

      //
      // --- support generating Extened VCD output by using
      //     '+define+tmax_vcde' on verilog compile line.
      //
      `ifdef tmax_vcde
         // extended VCD, see IEEE Verilog P1364.1-1999 Draft 2
         if (verbose >= 2) $display("// %t : opening Extended VCD output file", $time);
         $dumpports( dut, "sim_vcde.out");
      `endif

      //
      // --- IDDQ PLI initialization
      //     User may activite by using '+define+tmax_iddq' on verilog compile line.
      //     Or by defining `tmax_iddq in this file.
      //
      `ifdef tmax_iddq
         if (verbose >= 3) $display("// %t : Initializing IDDQ PLI", $time);
         $ssi_iddq("dut AAA_tmax_testbench_1_16.dut");
         $ssi_iddq("verb on");
         $ssi_iddq("cycle 0");
         //
         // --- User may select one of the following two methods for fault seeding:
         //     #1 faults seeded by PLI (default)
         //     #2 faults supplied in a file
         //     Comment out the unused lines as needed (precede with '//').
         //     Replace the 'FAULTLIST_FILE' string with the actual file pathname.
         //
         $ssi_iddq("seed SA AAA_tmax_testbench_1_16.dut");   // no file, faults seeded by PLI
         //
         // $ssi_iddq("scope AAA_tmax_testbench_1_16.dut");   // set scope for faults from a file
         // $ssi_iddq("read_tmax FAULTLIST_FILE"); // read faults from a file
         //
      `endif

      POnames[0] = "N387";
      POnames[1] = "N388";
      POnames[2] = "N478";
      POnames[3] = "N482";
      POnames[4] = "N484";
      POnames[5] = "N486";
      POnames[6] = "N489";
      POnames[7] = "N492";
      POnames[8] = "N501";
      POnames[9] = "N505";
      POnames[10] = "N507";
      POnames[11] = "N509";
      POnames[12] = "N511";
      POnames[13] = "N513";
      POnames[14] = "N515";
      POnames[15] = "N517";
      POnames[16] = "N519";
      POnames[17] = "N535";
      POnames[18] = "N537";
      POnames[19] = "N539";
      POnames[20] = "N541";
      POnames[21] = "N543";
      POnames[22] = "N545";
      POnames[23] = "N547";
      POnames[24] = "N549";
      POnames[25] = "N551";
      POnames[26] = "N553";
      POnames[27] = "N556";
      POnames[28] = "N559";
      POnames[29] = "N561";
      POnames[30] = "N563";
      POnames[31] = "N565";
      POnames[32] = "N567";
      POnames[33] = "N569";
      POnames[34] = "N571";
      POnames[35] = "N573";
      POnames[36] = "N582";
      POnames[37] = "N643";
      POnames[38] = "N707";
      POnames[39] = "N813";
      POnames[40] = "N881";
      POnames[41] = "N882";
      POnames[42] = "N883";
      POnames[43] = "N884";
      POnames[44] = "N885";
      POnames[45] = "N889";
      POnames[46] = "N945";
      POnames[47] = "N1110";
      POnames[48] = "N1111";
      POnames[49] = "N1112";
      POnames[50] = "N1113";
      POnames[51] = "N1114";
      POnames[52] = "N1489";
      POnames[53] = "N1490";
      POnames[54] = "N1781";
      POnames[55] = "N10025";
      POnames[56] = "N10101";
      POnames[57] = "N10102";
      POnames[58] = "N10103";
      POnames[59] = "N10104";
      POnames[60] = "N10109";
      POnames[61] = "N10110";
      POnames[62] = "N10111";
      POnames[63] = "N10112";
      POnames[64] = "N10350";
      POnames[65] = "N10351";
      POnames[66] = "N10352";
      POnames[67] = "N10353";
      POnames[68] = "N10574";
      POnames[69] = "N10575";
      POnames[70] = "N10576";
      POnames[71] = "N10628";
      POnames[72] = "N10632";
      POnames[73] = "N10641";
      POnames[74] = "N10704";
      POnames[75] = "N10706";
      POnames[76] = "N10711";
      POnames[77] = "N10712";
      POnames[78] = "N10713";
      POnames[79] = "N10714";
      POnames[80] = "N10715";
      POnames[81] = "N10716";
      POnames[82] = "N10717";
      POnames[83] = "N10718";
      POnames[84] = "N10729";
      POnames[85] = "N10759";
      POnames[86] = "N10760";
      POnames[87] = "N10761";
      POnames[88] = "N10762";
      POnames[89] = "N10763";
      POnames[90] = "N10827";
      POnames[91] = "N10837";
      POnames[92] = "N10838";
      POnames[93] = "N10839";
      POnames[94] = "N10840";
      POnames[95] = "N10868";
      POnames[96] = "N10869";
      POnames[97] = "N10870";
      POnames[98] = "N10871";
      POnames[99] = "N10905";
      POnames[100] = "N10906";
      POnames[101] = "N10907";
      POnames[102] = "N10908";
      POnames[103] = "N11333";
      POnames[104] = "N11334";
      POnames[105] = "N11340";
      POnames[106] = "N11342";
      POnames[107] = "N241_O";
      nofails = 0; pattern = -1; lastpattern = 0;
      prev_pat = -2; error_banner = -2;
      /*** No test setup procedure ***/


      /*** Non-scan test ***/

      if (verbose >= 1) $display("// %t : Begin patterns, first pattern = 0", $time);
pattern = 0; // 0
ALLPIS = 207'b011110000011001101110000100100111000110010110011011001111010100011101000101101100100101101001100010010100111101011100001110101011101000010101101100111000000001011001001110101110111111110001110011110000010101;
XPCT = 108'b000110101011111111000111001110000010011111111011011010001111010010011111000101101000110000011001001000111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 200

pattern = 1; // 200
ALLPIS = 207'b001111000001100110111000010010011100011001011001101100111101010001110100010110110010010110100110001001010011110101110000111010101110100001010110110011100000000101100100111010111011111111000111001111000001010;
XPCT = 108'b000111011101111111100011100111000001001111111001010000011111110011001111110101000010110000000001111001011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 400

pattern = 2; // 400
ALLPIS = 207'b011001100011111110101100101101110110111110011111101111100100001011010010100110111101100110011111010110001110010001011001101000001010010010000110111110110000001001111011101000101010000001101101111001100010000;
XPCT = 108'b001101001101000000110110111101100010110011111011111110011111101100010111011110001100111011111000111011111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 600

pattern = 3; // 600
ALLPIS = 207'b110010110010110010100110110010000011101101111100101110001000100110000001111110111010011110000011111001100000100011001101000001011000001011101110111000011000001111110100000001100010111110111000100010110011101;
XPCT = 108'b110000001001011111011100010010110011000011111101011011111111011110101111010101101111110000000000100010010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 800

pattern = 4; // 800
ALLPIS = 207'b000111011010010100100011111101111001000100001101001110111110110000101000010010111001100010001101101110010111111010000111010101110001000111011010111011001100001100110011110101000110100001010010001111011011011;
XPCT = 108'b001110100011010000101001000111011011010101101001011010010000100111111110110000100111101010111111111110111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1000

pattern = 5; // 1000
ALLPIS = 207'b100011101101001010010001111110111100100010000110100111011111011000010100001001011100110001000110110111001011111101000011101010111000100011101101011101100110000110011001111010100011010000101001000111101101101;
XPCT = 108'b110111011001101000010100100011101101010101111110001011001111000101101111000100001111110011011000110101010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1200

pattern = 6; // 1200
ALLPIS = 207'b101111110101101000111000011011100110100011110000001010010101001111100010101001001010110101101111001001000010010101000000000000000001010011011011001001110011001000000101001000100110010110011010111101110100011;
XPCT = 108'b110001001011001011001101011101110100010111111101011011011111000111111111101111000111110101111001010100101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1400

pattern = 7; // 1400
ALLPIS = 207'b010111111010110100011100001101110011010001111000000101001010100111110001010100100101011010110111100100100001001010100000000000000000101001101101100100111001100100000010100100010011001011001101011110111010001;
XPCT = 108'b001100100001100101100110101110111010001111111011011010011111011110111111101110000011111101100000110000001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1600

pattern = 8; // 1600
ALLPIS = 207'b010101111110010111111110100010000001011010001111011011011111110000010000000111110110000000010111100000110111001110110001110101011101010110011011010101011100111001001000100111111110011011101000110001011111101;
XPCT = 108'b000100111111001101110100011001011111101011111011111110001001010001111110000111100110111000000001011110111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1800

pattern = 9; // 1800
ALLPIS = 207'b001010111111001011111111010001000000101101000111101101101111111000001000000011111011000000001011110000011011100111011000111010101110101011001101101010101110011100100100010011111111001101110100011000101111110;
XPCT = 108'b000010011111100110111010001100101111001011111011011010011111101111111111011111001001110010000111001110001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2000

pattern = 10; // 2000
ALLPIS = 207'b100101011111100101111111101000100000010110100011110110110111111100000100000001111101100000000101111000001101110011101100011101010111010101100110110101010111001110010010001001111111100110111010001100010111111;
XPCT = 108'b111001001111110011011101000100010111101111111101111111001111011110110111011111011101111101111001100110010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2200

pattern = 11; // 2200
ALLPIS = 207'b101100101100111111001111010000101000111001100010100010100001011101101010101101011010011101001110101110100001010010010111111011110110101000011110111101101011101100000000110001001000001101010011011000001001010;
XPCT = 108'b110110000100000110101001101100001001100011111101111111110000101010100100011000111010100100011111100110100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2400

pattern = 12; // 2400
ALLPIS = 207'b101000010101010010010111001100101100101110000010001000101010001101011101111011001001100011101011000101110111000010101010001000100110010110100010111001110101111101001001101101010011111000100111110010000110000;
XPCT = 108'b110101100001111100010011111010000110111001111100101111011111100001011111100100100110111000111110011110001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2600

pattern = 13; // 2600
ALLPIS = 207'b110100001010101001001011100110010110010111000001000100010101000110101110111101100100110001110101100010111011100001010101000100010011001011010001011100111010111110100100110110101001111100010011111001000011000;
XPCT = 108'b110110111100111110001001111101000011100011111101111111001111111111101111010101001010110000100000101010100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2800

pattern = 14; // 2800
ALLPIS = 207'b100100000110011001010101010111110011111001010011111011110000000000111111110011010110110101110110100011111010011011001011010111010100100111000101001001011101010100011011101110100011000000000111100010100011001;
XPCT = 108'b111101111001100000000011110010100011110001111110100101011111111110001111001100110100111111100000101111110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3000

pattern = 15; // 3000
ALLPIS = 207'b010111000010101011100101110001000100001100100111100111000110100011100111010001010001000000010001111010011001001101010011000000101000001011011100110101010111011110001111001110011111001110001111100110101010011;
XPCT = 108'b001001110111100111000111110010101010011111111011011010010000000101101110000000010010101000000110000111011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3200

pattern = 16; // 3200
ALLPIS = 207'b010101100010011000000010011100011010110100100000101010011001110010011011000101001100001101000100101111101011001101001000010101001001000111000011111101101011100100001110010010111000011001001001101101010111100;
XPCT = 108'b001010011100001100100100110101010111101111111001111110001111000010001101110110100111111110100000010000111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3400

pattern = 17; // 3400
ALLPIS = 207'b101010110001001100000001001110001101011010010000010101001100111001001101100010100110000110100010010111110101100110100100001010100100100011100001111110110101110010000111001001011100001100100100110110101011110;
XPCT = 108'b111001000110000110010010011010101011011101111111011011001111110111001111100110110101110011111111000011111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3600

pattern = 18; // 3600
ALLPIS = 207'b101010101100010011000000010011100011010110100100000101010011001110010011011000101001100001101000100101111101011001101001000010101001001000111000011111101101011100100001110010010111000011001001001101101010111;
XPCT = 108'b110110010011100001100100100101101010011101111111011011010000000011001110101010111000101110111001101010001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3800

pattern = 19; // 3800
ALLPIS = 207'b010101010110001001100000001001110001101011010010000010101001100111001001101100010100110000110100010010111110101100110100100001010100100100011100001111110110101110010000111001001011100001100100100110110101011;
XPCT = 108'b000111000101110000110010010010110101100111111001111110010000010001101100000001110100101111011110010011000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4000

pattern = 20; // 4000
ALLPIS = 207'b010100101000001001000000100000000000000111011010011000101110010000001100011011101110110101010110011011111000111101111011100101110111010000100011100000111011011100000001101001010010001110111100001101011000000;
XPCT = 108'b000101000001000111011110000101011000111111111001111110011111010111111111000110000110110011100000000111101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4200

pattern = 21; // 4200
ALLPIS = 207'b010100010111001001010000110100111000110001011110010101101101101011101110100000010011110111100111011111011011110101011100000111100110101010111100010111011101100101001001000001011110111001010000011000101110101;
XPCT = 108'b000000000111011100101000001100101110111011111011111110011111111100101111101101011101111000011111010110010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4400

pattern = 22; // 4400
ALLPIS = 207'b010100001000101001011000111110100100101010011100010011001100010110011111111101101101010110111111111101001010010001001111110110101110010111110011101100101110111001101101010101011000100010100110010010010101111;
XPCT = 108'b000010100100010001010011001010010101111011111011111110010110000011011111100011011001101110011110001011001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4600

pattern = 23; // 4600
ALLPIS = 207'b001010000100010100101100011111010010010101001110001001100110001011001111111110110110101011011111111110100101001000100111111011010111001011111001110110010111011100110110101010101100010001010011001001001010111;
XPCT = 108'b001101011110001000101001100101001010000010111011011010010000110111111110111011000100101101111000010100110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4800

pattern = 24; // 4800
ALLPIS = 207'b111011000001000111100110101011010001111000010100011101001001100110001111010010111111111000100011101101110101001111110010001000110110100111010001011100001011100101010010100000100001110110100111111010100111110;
XPCT = 108'b111100001000111011010011111110100111000011110111011011101111110011101111111101101010110000111110110011100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5000

pattern = 25; // 5000
ALLPIS = 207'b111101100000100011110011010101101000111100001010001110100100110011000111101001011111111100010001110110111010100111111001000100011011010011101000101110000101110010101001010000010000111011010011111101010011111;
XPCT = 108'b110010000000011101101001111101010011111111111101111111100000000010000110101001101011101001111110011011000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5200

pattern = 26; // 5200
ALLPIS = 207'b100000110011011100001001001110001100101100110110011110101000111010001011011001001011010011000100101001111010111000011101010111010000101011011001110000000010110010011101011101111111100011100111100000101011010;
XPCT = 108'b110011101111110001110011110000101011111011111100101111001111010000111111000111100011111101111001011100010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5400

pattern = 27; // 5400
ALLPIS = 207'b110000011001101110000100100111000110010110011011001111010100011101000101101100100101101001100010010100111101011100001110101011101000010101101100111000000001011001001110101110111111110001110011110000010101101;
XPCT = 108'b111101111111111000111001111000010101101011111111111111101111100011101111011111000100111011011110101001001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5600

pattern = 28; // 5600
ALLPIS = 207'b111000001100110111000010010011100011001011001101100111101010001110100010110110010010110100110001001010011110101110000111010101110100001010110110011100000000101100100111010111011111111000111001111000001010110;
XPCT = 108'b111010110111111100011100111100001010111011111111111111010110001000001111001010011001100111000110100100100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5800

pattern = 29; // 5800
ALLPIS = 207'b111100000110011011100001001001110001100101100110110011110101000111010001011011001001011010011000100101001111010111000011101010111010000101011011001110000000010110010011101011101111111100011100111100000101011;
XPCT = 108'b111101011111111110001110011100000101110111111111111111110000100110100100000000110100100000000111001000111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6000

pattern = 30; // 6000
ALLPIS = 207'b101000111101000000001010010110011010100010101101011011000100110110000111101100010010101110110001011110001010010001111100001010111000010110001111111011110010111101111001011111010101100101101101100011101111011;
XPCT = 108'b110011110010110010110110110011101111111011111110101111101111000100001111100100000001110110100001100001000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6200

pattern = 31; // 6200
ALLPIS = 207'b110100011110100000000101001011001101010001010110101101100010011011000011110110001001010111011000101111000101001000111110000101011100001011000111111101111001011110111100101111101010110010110110110001110111101;
XPCT = 108'b110101111101011001011011011001110111100010111111111111011111100011011111010101010100111100000000111110011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6400

pattern = 32; // 6400
ALLPIS = 207'b110010110010010000001000110011111100001010000110001101110101111011100110010111010110000101011101001001101000110101100011001000010110010011101100000101001110010010100111001000100000111100110110111011010100101;
XPCT = 108'b111001001000011110011011011111010100010011011111011011001111101111011111001110010101110000000001010011011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6600

pattern = 33; // 6600
ALLPIS = 207'b110001100100001000001110001111100100100111101110011101111110001011110100100111111001101100011111111010111110001011001101101110110011011111111001111001010101110100101010111011000101111011110110111110000101001;
XPCT = 108'b111111010010111101111011011110000101100111111111111111111001100010011110101111100000110111100000111110101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6800

pattern = 34; // 6800
ALLPIS = 207'b010000001111000100001101010001101000110001011010010101111011110011111101111111101110011000111110100011010101010100011010111101100001111001110011000111011000000111101100000010110111011000010110111100101101111;
XPCT = 108'b000000011011101100001011011100101101101111111011111110001111011111011111011100011101111001100111101001100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7000

pattern = 35; // 7000
ALLPIS = 207'b101000000111100010000110101000110100011000101101001010111101111001111110111111110111001100011111010001101010101010001101011110110000111100111001100011101100000011110110000001011011101100001011011110010110111;
XPCT = 108'b111000000101110110000101101110010110101101111101110101111111010001101111110111111111110001111111011110010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7200

pattern = 36; // 7200
ALLPIS = 207'b011100111110110001001001000010000000101110111011111110011010001010111000110011101001001000111110110110111111000100111010100101100000001000010011001010000100111100000010011111111000010011101000001100100100000;
XPCT = 108'b001011111100001001110100000100100100101111111001111110010000100110101010010000110011101110111110010000100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7400

pattern = 37; // 7400
ALLPIS = 207'b101110011111011000100100100001000000010111011101111111001101000101011100011001110100100100011111011011011111100010011101010010110000000100001001100101000010011110000001001111111100001001110100000110010010000;
XPCT = 108'b110001111110000100111010000010010010011101111111011011001111111111001111101100010101111100111000001011110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7600

pattern = 38; // 7600
ALLPIS = 207'b011111110010101100011000000110111010101001000011100100100010010100101001100000101000111100111110110011100101100000110010100011100000010100001011001001010011110010111001111000101011100001010111100000100110011;
XPCT = 108'b000111001101110000101011110000100110010011111001011010010000011101111110000000110010101110111110101011000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7800

pattern = 39; // 7800
ALLPIS = 207'b010111111100101011000110000001101110101010010000111001001000100101001010011000001010001111001111101100111001011000001100101000111000000101000010110010010100111100101110011110001010111000010101111000001001100;
XPCT = 108'b001011110101011100001010111100001001000011111011011010000000001001011110110001010101101001111110001001000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8000

pattern = 40; // 8000
ALLPIS = 207'b000011000011010101101001010110101101110111100101000111100000100100100010100000010111101001010110101000010110111101111010011110100100010100101110100010111000100011101110010000010000111001100111011111101011101;
XPCT = 108'b001010000000011100110011101111101011001111101010001010001111101001101111010101101011111010111001010110010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8200

pattern = 41; // 8200
ALLPIS = 207'b101001011100101010111110111101001100011001011111111000110100100100010110111100011001011010011010001010000001001111000001000101101010011100011000101010101110101100001110010111011101111001011110001100011010101;
XPCT = 108'b111010110110111100101111000100011010101111111100101111100000111010001110111011011100101001011110010110110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8400

pattern = 42; // 8400
ALLPIS = 207'b100010101010001010100101111001001001100100111010100101001001111111000010000011010100111000010111111100101010000010001100011011100010110001001001110001011001010110111010111010100010111011111010000000101001110;
XPCT = 108'b111111011001011101111101000000101001000001111110001011110000110111011110011001000000101000111001000000011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8600

pattern = 43; // 8600
ALLPIS = 207'b110001010101000101010010111100100100110010011101010010100100111111100001000001101010011100001011111110010101000001000110001101110001011000100100111000101100101011011101011101010001011101111101000000010100111;
XPCT = 108'b110011100000101110111110100000010100111011111101111111101111110011111111101100010101111000100111111000000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8800

pattern = 44; // 8800
ALLPIS = 207'b010000110110110001011011110010011110111111011100100010001111100010111100001010000001011110101011001110101010001001010011101100111000001011000001001000000000101001110010100111101011000000000100000010011101111;
XPCT = 108'b001100111101100000000010000010011101100011111001111110010000011000101110111011111110101110000110111011110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9000

pattern = 45; // 9000
ALLPIS = 207'b001000011011011000101101111001001111011111101110010001000111110001011110000101000000101111010101100111010101000100101001110110011100000101100000100100000000010100111001010011110101100000000010000001001110111;
XPCT = 108'b000010011010110000000001000001001110111011111010101110001111001100001111101100101001111110100111000001000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9200

pattern = 46; // 9200
ALLPIS = 207'b000100001101101100010110111100100111101111110111001000100011111000101111000010100000010111101010110011101010100010010100111011001110000010110000010010000000001010011100101001111010110000000001000000100111011;
XPCT = 108'b000101001101011000000000100000100111101001111000101110001111000111101111011110010110111100011111001100010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9400

pattern = 47; // 9400
ALLPIS = 207'b100010000110110110001011011110010011110111111011100100010001111100010111100001010000001011110101011001110101010001001010011101100111000001011000001001000000000101001110010100111101011000000000100000010011101;
XPCT = 108'b111010101110101100000000010000010011001011111100001011111111000010001111111111111011111000100001100101011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9600

pattern = 48; // 9600
ALLPIS = 207'b010000011100101101101000100001111110011111010011100010000000101001000010010100000110101100001100001000010111000101101110101101100001100110011001111001100010111100101010111010011010110011101101101011101011100;
XPCT = 108'b001111010101011001110110110111101011101011111001111110001111111010101111111100100010111100100000100000111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9800

pattern = 49; // 9800
ALLPIS = 207'b100000110011010110111110000110100101101101000100101010000100100010100110100110010001111000110111011010000001110011001011011100001000100101000011000111000011100011101100000010011000111100011011010110011010101;
XPCT = 108'b110000010100011110001101101010011010101111111100101111101111100001111111110101111111110000011110111111110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10000

pattern = 50; // 10000
ALLPIS = 207'b011000100100101011010101010101001000010100001111001110000110100111010100111111011010010010101010110011001010101000011001100100111100000100101110011000010011001100001111011110011001111011100000001000100010001;
XPCT = 108'b001011110100111101110000000100100010111011111001111110011111101011110101001100000011111000000000101011001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10200

pattern = 51; // 10200
ALLPIS = 207'b101100010010010101101010101010100100001010000111100111000011010011101010011111101101001001010101011001100101010100001100110010011110000010010111001100001001100110000111101111001100111101110000000100010001000;
XPCT = 108'b111101110110011110111000000000010001110111111111111111100000011010111110100000000100100001011111000110010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10400

pattern = 52; // 10400
ALLPIS = 207'b011110110100001010111111000011001000100111101110101000100101011111110010100011100100001010011011110010111000111011111010010011110111010111000100011101110110001110111010101000110011111011010101100001100111111;
XPCT = 108'b001101001001111101101010110001100111001011111001011010010000101100001110110000110110101000111110111110010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10600

pattern = 53; // 10600
ALLPIS = 207'b001111010000000010100101100110101000101011010110110001001101100001111011000100101011101100010111100010100100011111000010101110000101100011111110111100101111011110010111110101011001011011011000111011110110100;
XPCT = 108'b001110100100101101101100011111110110011001111011010000000000100000010110101010011000101001111111101010000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10800

pattern = 54; // 10800
ALLPIS = 207'b000111101000000001010010110011010100010101101011011000100110110000111101100010010101110110001011110001010010001111100001010111000010110001111111011110010111101111001011111010101100101101101100011101111011010;
XPCT = 108'b001111011110010110110110001101111011010101111000000000010000000101101100011000101001101100000110000000001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11000

pattern = 55; // 11000
ALLPIS = 207'b100011110100000000101001011001101010001010110101101100010011011000011110110001001010111011000101111000101001000111110000101011100001011000111111101111001011110111100101111101010110010110110110001110111101101;
XPCT = 108'b110111100011001011011011000110111101011111110101011011100000110011011110101000110101101010011110010001101001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11200

pattern = 56; // 11200
ALLPIS = 207'b100110100101010000111010110010100111010100010011100011010011100101000101110101001110001111110111001010100000110001000101010100010111101011001001110000110101010001001001010001111001110111100010011001000001011;
XPCT = 108'b110010001100111011110001001101000001011011111110001011101111101011001111100100011001110100111111101100101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11400

pattern = 57; // 11400
ALLPIS = 207'b100001010110111101111111001110000000000101100000001101111111110110100110000001010101100001101000010010000101110011011001000101100111010110010000000111011110111100101111000011110111111101110011111000100001100;
XPCT = 108'b111000011011111110111001111100100001111011111110101111001111100111000111001101100110110101100000010100011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11600

pattern = 58; // 11600
ALLPIS = 207'b100010101111001011011101110000010011101101011001111010101001111111010111111011011000010110100111111110010111010010010111001101011111001000111100111100101011001010011100001010110000111000111011001000010001111;
XPCT = 108'b110001011000011100011101100100010001001011111100001011001111011001001111111110100111111000100110111101110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11800

pattern = 59; // 11800
ALLPIS = 207'b110001010111100101101110111000001001110110101100111101010100111111101011111101101100001011010011111111001011101001001011100110101111100100011110011110010101100101001110000101011000011100011101100100001000111;
XPCT = 108'b111000100100001110001110110000001000101111111111111111101111011111111111001110111111111000100111101100010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12000

pattern = 60; // 12000
ALLPIS = 207'b010101010111110011101010100101101011101010011111110001011110001101111000100010100010010001111101000100011000001111101111001110011101101000111101111000000111010011010110010100110011100100000110000011000010101;
XPCT = 108'b001010101001110010000011000011000010101011110011111110001111101110111111111101011101110000111000101001100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12200

pattern = 61; // 12200
ALLPIS = 207'b011000101111101100010111000101100110011010100110000100111001000010111000101010100011101110101101010101011001101100001100001000100010010111101010000011000111111101100000100001010010110100000001110101100000011;
XPCT = 108'b000100000001011010000000111001100000101111111001111110001111010111000101011110001110110100011110001111111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12400

pattern = 62; // 12400
ALLPIS = 207'b001001000001101000000000101111111111011100111101001100110001001100010011111110100110111011100110011101111110100110011010001110101000110001001001101111011100101011100111101111000001010000100010111010101101001;
XPCT = 108'b001101110000101000010001011110101101110001111001111110011111100101011111000111101011110111011001010101111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12600

pattern = 63; // 12600
ALLPIS = 207'b110110100100100001100010000000101100000001110111011010001110100010001101000100100001111011100000111001101010111000110110101000111000111011010000001000101010000001111000011100101011101110010011101001010111101;
XPCT = 108'b110011101101110111001001110101010111000011111101011011111111101010111111110100010011110010100001000001100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12800

pattern = 64; // 12800
ALLPIS = 207'b001111101101011101111010110111011000101111110100001010110101101100100111101010111010111000101011111001001111000101110110000101100010101101000000111101001110110100010101101100000001111101100110001110010100110;
XPCT = 108'b000101100000111110110011000110010100010111111001011010001111101110010111101110100110110000100110011000100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13000

pattern = 65; // 13000
ALLPIS = 207'b110001111111000010111100111010100101100100010100111110111011011111001101000001011100001000011001001001000110011010100110001110110100001000100100110000010111111001001110110000001011011001011011010111100100000;
XPCT = 108'b111110000101101100101101101011100100100111111101111111111111001001001111011111111100111110111001000000001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13200

pattern = 66; // 13200
ALLPIS = 207'b100101011101111010011110000101000000101110110001110001100101110101110001001101101110010001001111101001111011010011010100010100011011010011110011010011100111110100010110011001100111010101010111101111111001100;
XPCT = 108'b111011001011101010101011110111111001100111111111110101001111101001111111111100000000111100111110011001100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13400

pattern = 67; // 13400
ALLPIS = 207'b110010101110111101001111000010100000010111011000111000110010111010111000100110110111001000100111110100111101101001101010001010001101101001111001101001110011111010001011001100110011101010101011110111111100110;
XPCT = 108'b111001101001110101010101111011111100011111111101011011110000000000110100000000000111101010111111111001110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13600

pattern = 68; // 13600
ALLPIS = 207'b111100101011101111010011110000101000000101110110001110001100101110101110001001101101110010001001111101001111011010011010100010100011011010011110011010011100111110100010110011001100111010101010111101111111001;
XPCT = 108'b111110010110011101010101011101111111100111111101111111001111100000011111111100011010111001111001110010111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13800

pattern = 69; // 13800
ALLPIS = 207'b001100010001100010001011101111000111101101010010111011010000010011010011111111000100011111010111001001110010000110110110111110111101001110111011110010001010001011011010110010101101011011010111101010111110101;
XPCT = 108'b001110011110101101101011110110111110100011110010101110001111000011001111110101111000111001011000110000010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14000

pattern = 70; // 14000
ALLPIS = 207'b111000000010000111110001100111001011100011001001101100101001000010110010011001111010110010101111111110100011111111101011110111110101100001100000011100000100111100111000110010000101110011110110010100101110000;
XPCT = 108'b110110010010111001111011001000101110100111111101111111001111010000001111011111101010111011100001100010110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14200

pattern = 71; // 14200
ALLPIS = 207'b111100000001000011111000110011100101110001100100110110010100100001011001001100111101011001010111111111010001111111110101111011111010110000110000001110000010011110011100011001000010111001111011001010010111000;
XPCT = 108'b110011000001011100111101100110010111100011110101111111101111000001101111111100010011111001011001001100111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14400

pattern = 72; // 14400
ALLPIS = 207'b001100000100110100011110001110100001010111011011100111011100010100101000011101101100001010111000001000111101010100000001010010010001111011101100111000000101011011000101100111101010011010111111010001001010101;
XPCT = 108'b000100111101001101011111101001001010110011011011111110010000100100000100000011111100101001111111110000011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14600

pattern = 73; // 14600
ALLPIS = 207'b100110000010011010001111000111010000101011101101110011101110001010010100001110110110000101011100000100011110101010000000101001001000111101110110011100000010101101100010110011110101001101011111101000100101010;
XPCT = 108'b111110011010100110101111110100100101001011111111011011000000100110101110010011101000100010111001001111110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14800

pattern = 74; // 14800
ALLPIS = 207'b010000100010101100010010111010011101111101001111100010110000100000100111011110010100110010011110111010101101011111011101111101100100011110100111111000100010100001011101011001011000110000010110100000001001110;
XPCT = 108'b000011000100011000001011010000001001111011111001111110011111001010111111001110010011111100100000111110011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15000

pattern = 75; // 15000
ALLPIS = 207'b111001011111111110000110011101111001101101011011010101110100010100100111000110111000110110100011100100111000110011100110111101010001101000101000011011010010001110000110011101110011100010111101100011101100110;
XPCT = 108'b111011101001110001011110110011101100101011111111111111001111111100011011011110110100111001100110100111000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15200

pattern = 76; // 15200
ALLPIS = 207'b000101110111111101101011000001010100101100111011001011000001111000100000111010100111010110001100010100000111011000010010101000100110100011110010101011000010110001101011000001001000011111101001111100001110010;
XPCT = 108'b001000000100001111110100111100001110110111111010101110011111101111001111110101101100111100011111010001100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15400

pattern = 77; // 15400
ALLPIS = 207'b001110111110111100100010101101000101001001111100011000001010101100011001101001111001001100100111011001001101000101111100110001001111010001011010101110010101001101000010101101010111110111011000111001001110000;
XPCT = 108'b001101100011111011101100011101001110001001111001011010010000000010001010011010000110100100111111100100010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15600

pattern = 78; // 15600
ALLPIS = 207'b000111011111011110010001010110100010100100111110001100000101010110001100110100111100100110010011101100100110100010111110011000100111101000101101010111001010100110100001010110101011111011101100011100100111000;
XPCT = 108'b000010111101111101110110001100100111010101111001011010011111100000011111110111101101111011011000011011100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15800

pattern = 79; // 15800
ALLPIS = 207'b010001010000010011000100010000100010001000101001101101101010000010001000010111101111111110001110111111100010110110010010110110110000100101000110011101000001001111011100010000110010111000001101001001001010001;
XPCT = 108'b000010001001011100000110100101001010101011111011111110010000001000101110111010101110100111011111011010011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16000

pattern = 80; // 16000
ALLPIS = 207'b110100010100000100110001000100001000100010001010011011011010100000100010000101111011111111100011101111111000101101100100101101101100001001010001100111010000010011110111000100001100101110000011010010010010100;
XPCT = 108'b111000100110010111000001101010010010110011110111111111101111101001011111000101011101110010100001001000100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16200

pattern = 81; // 16200
ALLPIS = 207'b100011010110101100111101010110000001010101000101011101100010001100010110010111010100010100000000001100011100010000110001011001101001001111101011111011100100111001100001001110010010111110110010100011011101110;
XPCT = 108'b110001110001011111011001010011011101011011111111011011000000011011101110100011110011101101000110000010010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16400

pattern = 82; // 16400
ALLPIS = 207'b010001101011010110011110101011000000101010100010101110110001000110001011001011101010001010000000000110001110001000011000101100110100100111110101111101110010011100110000100111001001011111011001010001101110111;
XPCT = 108'b000100110100101111101100101001101110100011111001111110001111011011111111110100011110110000100000110000011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16600

pattern = 83; // 16600
ALLPIS = 207'b011010001010010111000011101110010011001111100111111100110000001010001011101000000100101000000111001010110110100011000001101100111001000010101010001000011101010010010100101000000011101010010111101111101110110;
XPCT = 108'b000101000001110101001011110111101110000111111001011010001001011100101110010100100110111010100001111110100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16800

pattern = 84; // 16800
ALLPIS = 207'b111111111101011011110110100110011101011110100010101010111000010110000101111100111001111100100010010110010101011011010110100110011111111000000010111001010101011010100011010111110011011000011000011000010111011;
XPCT = 108'b111010111001101100001100001100010111011011111101011011110110001111010111100001001011101001111110000110110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17000

pattern = 85; // 17000
ALLPIS = 207'b011111111110101101111011010011001110101111010001010101011100001011000010111110011100111110010001001011001010101101101011010011001111111100000001011100101010101101010001101011111001101100001100001100001011101;
XPCT = 108'b000101011100110110000110000100001011011111111011011010000000000110101110100010100100100010111111011100010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17200

pattern = 86; // 17200
ALLPIS = 207'b011011110000000000010010011110010000011100011110110110001100001111101100101101101001111001001001111101000011011000000011001111111100010010010100100010100110000000010011001011111010100101000000001101011011010;
XPCT = 108'b001001011101010010100000000101011011011111011001011010010000111101111110100000110000101101111000111010010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17400

pattern = 87; // 17400
ALLPIS = 207'b001101111000000000001001001111001000001110001111011011000110000111110110010110110100111100100100111110100001101100000001100111111110001001001010010001010011000000001001100101111101010010100000000110101101101;
XPCT = 108'b000100101110101001010000000010101101111111111010100100000000111110111110000010001100101101011111100110111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17600

pattern = 88; // 17600
ALLPIS = 207'b111010000001111110000100001110001011101110111000100011000101110101011010100011010101111001101010101011010000101000100110100100101110001010111010111111000110111110000100000100101100110110010101100010000111101;
XPCT = 108'b110000101110011011001010110010000111000011111111011011111111111011101111010110011101110100011110111011001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17800

pattern = 89; // 17800
ALLPIS = 207'b101111111111000011001110111100110110101101101010111010001010010011100011011100011011010001110010011100011001110011011110101000110100010100001101101001000111000011001110111001110001011110110001110110011010011;
XPCT = 108'b111111001000101111011000111010011010001111011100001011011111111111011101011110110010110001111001111000010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18000

pattern = 90; // 18000
ALLPIS = 207'b100101111111111000011001110111100110110101101101010111010001010010011100011011100011011010001110010011100011001110011011110101000110100010100001101101001000111000011001110111001110001011110110001110110011010;
XPCT = 108'b110110110111000101111011000110110011110111111110101111111111110000011101000111000011111001100001111100111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18200

pattern = 91; // 18200
ALLPIS = 207'b011100100110111101010000100001001110101001010000111101101011110110111111111010011010001011010001010101110010100100000111110101000110111011001100110100001010110101101101000001110110010010110101010111000110010;
XPCT = 108'b000000001011001001011010101011000110111111111011111110000000100100111010001000011101101110011111000100110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18400

pattern = 92; // 18400
ALLPIS = 207'b001100011001110110110100001101101000110100111111101111110010101000100100010000101110100001101100000010111101011010111100011000101011101111000000100101011110001101000011110100110010001010101010000100000110111;
XPCT = 108'b001110101001000101010101000000000110111101111011111110011001011001111110100111001000111011100110100011011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18600

pattern = 93; // 18600
ALLPIS = 207'b100110001100111011011010000110110100011010011111110111111001010100010010001000010111010000110110000001011110101101011110001100010101110111100000010010101111000110100001111010011001000101010101000010000011011;
XPCT = 108'b110111010100100010101010100010000011011011111111011011010000111010011110000011100000100110111001001011000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18800

pattern = 94; // 18800
ALLPIS = 207'b010011000110011101101101000011011010001101001111111011111100101010001001000100001011101000011011000000101111010110101111000110001010111011110000001001010111100011010000111101001100100010101010100001000001101;
XPCT = 108'b000111100110010001010101010001000001000011111011011010001001111010001110101101110000111111000000111100011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19000

pattern = 95; // 19000
ALLPIS = 207'b000110110001010101011100100000110101100111100111001100001000000111011101000000110010000010110011011011010101101110000100100111000010010100100010010100100011001010110011100000110100101100111011101001110010001;
XPCT = 108'b001100001010010110011101110101110010011011111001011010011111111001111111000111001110110010011110011111100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19200

pattern = 96; // 19200
ALLPIS = 207'b100100010000110111111011000101001000000101101100000100001010110110000100010010011100011011000111001110101000001001110111010001111110101001101000100110101110101100111011011101110000110111010010001010001000000;
XPCT = 108'b111011101000011011101001000110001000111011111100101111111111111111001011100110000011110100100001111101001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19400

pattern = 97; // 19400
ALLPIS = 207'b001110001100101000010000001100101110111000100110100100110110000110110010111000111111110111011100101111101011000011011010001110000101101100011101001110011100101001101000101101011010110010110001111010010101010;
XPCT = 108'b000101100101011001011000111110010101001001111000000000000000111011111110110010100110101100111001110011101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19600

pattern = 98; // 19600
ALLPIS = 207'b100111000110010100001000000110010111011100010011010010011011000011011001011100011111111011101110010111110101100001101101000111000010110110001110100111001110010100110100010110101101011001011000111101001010101;
XPCT = 108'b110010111110101100101100011101001010000111011101011011101111111011001111101101000100111011100000100010100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19800

pattern = 99; // 19800
ALLPIS = 207'b100011101010101001001011000001101010011010100010101011100101001010000010101001010100001001100011001001111100101001011110101100111111011111101011100100110001001001111101011100100111010110100101111110111011101;
XPCT = 108'b110011101011101011010010111110111011010111111110001011100000000001101110100001101111101010111110110000001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20000

pattern = 100; // 20000
ALLPIS = 207'b110111101001000010010100101110100001100010011001011000100101101000000010011110010100110010100000010111000110100011000100001011101010111111111100100100001100011011001000110101111011001100000001011011111011110;
XPCT = 108'b110110101101100110000000101111111011001011011101011011001111101101110111100101101010111100011000101010000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20200

pattern = 101; // 20200
ALLPIS = 207'b111010010011011101010000001011000100001000000110001110110010010011001100010110111110110111110111011000010000101010011000100000111001001011010010000001000111011011011111110010010111101101110111001010010111100;
XPCT = 108'b111110010011110110111011100110010111011011111101011011011111111001111011000111101010110001111110000111111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20400

pattern = 102; // 20400
ALLPIS = 207'b101110101010000000001101111010000111001001100101010110010011010001000110110010001001011100110011101111110100000101010111100110000011111011101001101001111110111001100100110011101000010100010110001100010011100;
XPCT = 108'b110110011100001010001011000100010011000111111101011011100000001110000100011000001010100110011111010010010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20600

pattern = 103; // 20600
ALLPIS = 207'b101110011100011110101100011100000111000001100010001111011110011100110111110010011101111101101101101110011000000000101001000011011011110000010001010010100111101111100011011001010000010000100000011101000000010;
XPCT = 108'b111011000000001000010000001101000000011111111111010001110000100101001110000000110001101110011111011011000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20800

pattern = 104; // 20800
ALLPIS = 207'b110111001110001111010110001110000011100000110001000111101111001110011011111001001110111110110110110111001100000000010100100001101101111000001000101001010011110111110001101100101000001000010000001110100000001;
XPCT = 108'b110101101100000100001000000110100000010111111111011011110000010011111100101011010101100000011110100001011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21000

pattern = 105; // 21000
ALLPIS = 207'b011000011001101011011101000011001001011101011111010000011111000100110011110101101010000100110011111111101011011111111101111000111110001010001110111000011110101100000010010011011101101010011100100001101000110;
XPCT = 108'b001010010110110101001110010001101000101011111001111110011111010111111111010111111011111001100110011011110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21200

pattern = 106; // 21200
ALLPIS = 207'b001111010010010010110101100010001000011011011101101100101010110000000000101010111010000101101111101001110010111010101000100101101001001001001000111010000101100011110010000101100000001000011001001010110110111;
XPCT = 108'b001000101000000100001100100110110110000001111001011010000000110100111110011000101111101100111001101110001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21400

pattern = 107; // 21400
ALLPIS = 207'b100111010100000111100110100101011111011001000011010011011110101101111111000110100111011110011101001101000001101011101001011101111101001011101000111100000000001110100000110111011011010010100011001000001001010;
XPCT = 108'b110110110101101001010001100100001001001001111111010001110000110011011110001010010111100111000111100101001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21600

pattern = 108; // 21600
ALLPIS = 207'b101001101110100011010111110001000011010010100110011011100011101000011010100111111101110100100111101111100100000001100000001000101010011111101100001001001111010010000000011111000011010001000011110101010110110;
XPCT = 108'b110011110001101000100001111001010110100101011111111111000000001011101010100000000000101101100111110100110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21800

pattern = 109; // 21800
ALLPIS = 207'b000110111101001110110110000111011001101011100100001001001010100100110010100000011110001111101100101100001110101010101100110011101100011000011111001100010101101011100110011000011101111010101110110100000101001;
XPCT = 108'b001011000110111101010111011000000101001101111011010000011111100101101111011111010001110111011111000010011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22000

pattern = 110; // 22000
ALLPIS = 207'b000111111100101011010001001000010000101110010100100000001010000110111000001001110110001001100000010010111010100001011100100101010000101101100101110100001110101110110000111000110000011001010011010101001000011;
XPCT = 108'b000111001000001100101001101001001000001101111001010000010000101111111110011001101001100001011110001011000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22200

pattern = 111; // 22200
ALLPIS = 207'b011011110010101000101100101000101100100100011100000011010011110110011000001000011010111101110000110001000111010000000110010100011000000001010110101000010100001011000101000000010011101010010110101110100000100;
XPCT = 108'b000000000001110101001011010110100000011111111011011010001111000110111111001111100010111011000000010101010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22400

pattern = 112; // 22400
ALLPIS = 207'b110001101100001110110000011100010110100000011011001010011011101110010000011100010011111110100100111011111011101000101010100110101011010110111010000011011010010001101100101001111011001000100100111000010100111;
XPCT = 108'b110101001101100100010010011100010100101011111101111111101001100011001110011101100001111100000001011010111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22600

pattern = 113; // 22600
ALLPIS = 207'b110111001000010101101100000101101001111110110111100100100100100001110010100100101110001011100011100010011000111010101101001100010110001110110111100110010000011010101101111110011110001001000111101100101101101;
XPCT = 108'b110111110111000100100011110100101101011111111101011011100000001010101110100001101101101110011110001001110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22800

pattern = 114; // 22800
ALLPIS = 207'b111011100100001010110110000010110100111111011011110010010010010000111001010010010111000101110001110001001100011101010110100110001011000111011011110011001000001101010110111111001111000100100011110110010110110;
XPCT = 108'b111111110111100010010001111010010110000111111101011011000110110000011111000010000000100000100111001100000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23000

pattern = 115; // 23000
ALLPIS = 207'b111111101111000011100110100100111100011110011010011100100111110001110101000100011100110011101010000101010100110110011010101010011011011010101101110101101111110000000101001010011111011110110111100110100101101;
XPCT = 108'b110001010111101111011011110010100101011111011101011011001111010101111101000101000111110001011000000110111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23200

pattern = 116; // 23200
ALLPIS = 207'b110100001000000000011101110101001100101010111100000000100010100110100000001101100101100111011100010000101110000110000000010111100010000101001001001111111110010101011010011111111100011011001011100101001010001;
XPCT = 108'b111011111110001101100101110001001010101111111101111111001111110011101111111101000011111001000001101001010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23400

pattern = 117; // 23400
ALLPIS = 207'b110001011010000000100001000010000110110101101011000001101111000010001000010101110111110000010011110101111001101011100000111101011110101110001001000011111101011010111000000111111011101011101110010110001100111;
XPCT = 108'b110000111101110101110111001010001100101110111111111111000000110110111110111010010110100001100110001000111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23600

pattern = 118; // 23600
ALLPIS = 207'b100011010111110100110111111100010010101000011010110111010011010100100000001100111110111110001101101100100101001100100111100111110011100101000011100011111011101000000111010011110110101111111100111000110100011;
XPCT = 108'b111010011011010111111110011100110100011001111111011011111111100000011111010110001101110110000000111101101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23800

pattern = 119; // 23800
ALLPIS = 207'b001100001010111110011101010101111011000000111011010111111111010111100100011010101100111001001001001100111000100101100100010011111010010110111010000011100011110111110100000101100110000011101000101101010010110;
XPCT = 108'b000000101011000001110100010101010010100111111011111110000000010010111110011010111101101111011000000100100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24000

pattern = 120; // 24000
ALLPIS = 207'b101110101101010101001010000100111101010011110000010111111111110100001011010100100000001000011111011001010111001110111011101110101110101100110010000101111011010101011101001011110010010100101100110101000010100;
XPCT = 108'b110001011001001010010110011001000010011110111110001011101111000000001111100100010101110110011000000001010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24200

pattern = 121; // 24200
ALLPIS = 207'b000010000000000111011101010011001010101111000000001000101001101000000011011001011001110111000100001011100001100000000101111000100001010010010011111111100101010110100111111111000110110010111001010010100010001;
XPCT = 108'b001111110011011001011100101010100010010011111001011010011111100001011111001101000010111100100001111011100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24400

pattern = 122; // 24400
ALLPIS = 207'b101111111100100000100110001000001110110101111100111000000011000100000111100000000010110001001011101010010110100000110001000011110111111111100011101011000010000000011011000010100111111011000001001110010100010;
XPCT = 108'b111000011011111101100000100110010100010101111100001011010000111101011010001001001111101000100110001110010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24600

pattern = 123; // 24600
ALLPIS = 207'b001011101100011101000101100110011110001001111100001110000101010010101011111100111110000100011100111110000010011111100101100000111111000101010000110010001010110111110110101100001111110100011011010101100111110;
XPCT = 108'b001101100111111010001101101001100111000101111001011010000000000100001110010011111011100111111001011010000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24800

pattern = 124; // 24800
ALLPIS = 207'b111101100000010110110111100000000001100011100100100101110001011001111000001001111100110101100100010010010100001001001001110001001101011111100000010000100001110110111000110000001110110101110010100100000101001;
XPCT = 108'b110110000111011010111001010000000101100111111111111111010000001000101100010011011000100100111111111011011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25000

pattern = 125; // 25000
ALLPIS = 207'b000011101000101111101010001101011000100011110110000011110101000110011000000010011101011001010000110011001000111101010011001010000000011011010001110010100000011101110010001110000101110001011101110001010001000;
XPCT = 108'b001001110010111000101110111001010001000011111011011010011111111000101111100100100011110110100000111111011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25200

pattern = 126; // 25200
ALLPIS = 207'b110011000010101000011111010101100011101100111100101010100101000000011000000000001001010000100111011110110111111100000101011001001100110010100111011010100000000001110000001000011001110000000101100001000001000;
XPCT = 108'b110001000100111000000010110001000001001011100101011011011001100010011110100111110010111100100000111010100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25400

pattern = 127; // 25400
ALLPIS = 207'b011001100001010100001111101010110001110110011110010101010010100000001100000000000100101000010011101111011011111110000010101100100110011001010011101101010000000000111000000100001100111000000010110000100000100;
XPCT = 108'b000000100110011100000001011000100000100011111011111110001111000000111111011100010010111001111111000111001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25600

pattern = 128; // 25600
ALLPIS = 207'b000111011110111101010101110001110101011010001101101000110101110101000001011110111110111101100001010011100111001111011101000110100010010000001011110001010100010101110101000001001001100010101010001000010111010;
XPCT = 108'b000000000100110001010101000100010111010000111001011010010110111111111111110001011111101010011111001000000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25800

pattern = 129; // 25800
ALLPIS = 207'b110000101100100101111011111011110010101111011000111100100001101101100000101001110011000011000111010010001110110000011010000100000010001010111110001011110101000100010110101100001111011101100110110110000110101;
XPCT = 108'b111101100111101110110011011010000110100111101101111111001111110011111111111110010110110000000000101100000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26000

pattern = 130; // 26000
ALLPIS = 207'b111011011110001001001110010000101101001100110000011010100110100100011010110001100001100010110010101001010011110110010000110010111101011100001011000111101111000001110101011100110101100100111100001111111110000;
XPCT = 108'b110011101010110010011110000111111110011111111101011011010000000110111100101001100011101100011111000010001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26200

pattern = 131; // 26200
ALLPIS = 207'b101011101110101011000111001010001000001011110010110010011101001010000000010011011001000010110010100111011001010001010001001010001111010111110101111111010100010100100010101010110011110101100111100111101111000;
XPCT = 108'b111101011001111010110011110011101111001101111101011011011001101010010100000111000110110001000000111100001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26400

pattern = 132; // 26400
ALLPIS = 207'b101110111111001111111010101111000001011010100101111101000000010111000011010011110111011001010011001001110111010000110100111010010111100001101010100100010111100110100001110000101100011001001101010111111011010;
XPCT = 108'b110110001110001100100110101011111011010111111111011011101001101001001010001111111000111001011001100000111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26600

pattern = 133; // 26600
ALLPIS = 207'b011011110101101111100000110010100111101110100111000001101010000111111111110111000101010001011001011101111110000101001100000110000001101000110000110000010000111101000111100100001111011000110001101111111001010;
XPCT = 108'b001100100111101100011000110111111001010111111011011010011111100111011101100101010000110101011000000100100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26800

pattern = 134; // 26800
ALLPIS = 207'b001100011101010011000010111100001010010100010001011110111111011100001110111101110111110100101000101011011111010000100011100111111001110010000001010001111100011001001101011011101110100000000100101101011001111;
XPCT = 108'b000011011111010000000010010101011001110101111000101110001111001110001111000111100011111110000001101100011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27000

pattern = 135; // 27000
ALLPIS = 207'b011111110010110110011001001001010010111000000110011100101000000110100011100101100011110110100001111000001111011101100111011001011101100011001110001001110101000100000110000111101010010110101101111101100101000;
XPCT = 108'b001000111101001011010110111101100101000111110001011010010000011001011110110011011111100101111110010111010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27200

pattern = 136; // 27200
ALLPIS = 207'b110001111010010011001101100100101000000110111001010111011111101010010010010110111100001001101010101100011110100011000111000010000010101111000010000101100011110101010110111011111101111011110100001101111100000;
XPCT = 108'b111111011110111101111010000101111100101111111111111111110000100111101110111000001101100100111110110010011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27400

pattern = 137; // 27400
ALLPIS = 207'b110010110001011101100101100111001110111001110000010011000000001001000000001111011011100111010111100011010011101110100011101101000000111000111111000000001001111010111010100010010001001100001001010100001011011;
XPCT = 108'b111100010000100110000100101000001011001111111111011011011111100101110101011111111100110010000111101111101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27600

pattern = 138; // 27600
ALLPIS = 207'b001001001001100000111001110111101011010000011000101100000110111000110000111011010000101000111011101101011001010000011010000111111011110001010110111010111100101000100001111010111111001111101000111001011010101;
XPCT = 108'b000111011111100111110100011101011010111011111001110100001111001101101111000100011000110000111001111010101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27800

pattern = 139; // 27800
ALLPIS = 207'b110011111000111111110000101110101111100100011101100111101111010001001001110110110000011001101011011011000001101011101101010101000010110100011101000010010110010001000001010100111010001101011111010110010011110;
XPCT = 108'b110010101101000110101111101010010011011111011111011011100000001111010110011010101010101110111001000011101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28000

pattern = 140; // 28000
ALLPIS = 207'b110111100101100111000010011110111001010001010111011001000101000111101100111001110100110001100111110011111010000001011011101111000111100000011101000000101000111100011010100011101100010111110100101011111101101;
XPCT = 108'b111100011110001011111010010111111101000011111111011011001111000111111111000100011110111101011000001100011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28200

pattern = 141; // 28200
ALLPIS = 207'b001001000110011001001101010010001010101110000000011000100100011010111111110111110111011000101101111110000011001011011100000000000000110011111100000101101011010110000111110101000100100101110110111100011100110;
XPCT = 108'b001110100010010010111011011100011100110111111001110100000110101111111011101001001010100110111111100110011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28400

pattern = 142; // 28400
ALLPIS = 207'b101011101001111011101110010101101111110001011001111110110110111000011101110100011110101010001111100001011011001110001011101001111001101000101101110110110001001110100101010000100011000000111001111000001110011;
XPCT = 108'b110010001001100000011100111100001110010011111101011011111111011001100111001100101110110001011000110000011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28600

pattern = 143; // 28600
ALLPIS = 207'b001110011111011001011100101011100010100001010111101010001011001011111011110100111110111111000111100010010000100110101010011011001100001101001000010001011001101110000101101011101001000100110000100001011001001;
XPCT = 108'b000101011100100010011000010001011001010011110001010000011111011111111111100111010110110111111000010001000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28800

pattern = 144; // 28800
ALLPIS = 207'b100001100101111101111000001001111000000100011110100101111011110101101010001010100011101010101011111001111110000111101110010111100000011011110000011000001000011110110101011010001001000100110011111000100111010;
XPCT = 108'b110011010100100010011001111100100111110011111111111111111111101000101111011110100000110001100110011001101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29000

pattern = 145; // 29000
ALLPIS = 207'b000001100111011011100100011001110100100001100101101010000110110100010000101110101111101100111100110100000100010111011101101100001110100010001100110111000110000000011000100110111111111011010000010111101011110;
XPCT = 108'b000100111111111101101000001011101011101101111000101110001111111011111111111111110111110010100001111010111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29200

pattern = 146; // 29200
ALLPIS = 207'b100011000010001100010111001110111101101100000000110000111001011011101100110111101101110000001001011010010101101111001000110101110111010001101111010001011101110001010100110111010110001001010111000000001011110;
XPCT = 108'b110110110011000100101011100000001011001000011101011011000000011100111110100001100001101010100110001000001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29400

pattern = 147; // 29400
ALLPIS = 207'b100011100001101111100000111111111011100011011110100111111011110001011010000001011010000101010000110110000111001101000101110001100000111110000000111110000011111011010011001100100011110100000001011000111011111;
XPCT = 108'b111001101001111010000000101100111011010001111111011011001111101101011111110111011101111001000110010011010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29600

pattern = 148; // 29600
ALLPIS = 207'b111101100100010011101001110001110111101001010010101110000000110000000011110101110101001001110001111011000110111110011000111000010111110111001111001110100110110010110110101001101010010111100001010111010100000;
XPCT = 108'b111101001101001011110000101011010100100111001101111111110000000000011000011000000110100110011110011101010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29800

pattern = 149; // 29800
ALLPIS = 207'b100111011010000000010011101101010010000111000000001000000110111001110011011010100100010011001101011100111000111011001010001010001001111100101110110111001111010101110100011010110010100011101100101100010001100;
XPCT = 108'b110011011001010001110110010100010001001101111101010001000000100010001110011000000110101001011111111001010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30000

pattern = 150; // 30000
ALLPIS = 207'b101011000101101110100110101001100011010100100101110110001010001001101110011100100101100001110001111010000100101100100001010101010011101101100011111110000000010110011111001111011010111101000111111000101110000;
XPCT = 108'b111001110101011110100011111100101110011001111100001011011111110100010111010100001101110011111001001100010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30200

pattern = 151; // 30200
ALLPIS = 207'b101100101100111111001110011100011001011011011011000110000110010001100100011010001111101111000000110001111110000101001101111101011110000001011011010100111110100010101010011001101000101000100101000100100010100;
XPCT = 108'b111011001100010100010010100000100010100111111100101111110000010001111110010000000011101011011110100001000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30400

pattern = 152; // 30400
ALLPIS = 207'b001101110010101110001001011101010100111101100100111101111010111011001010000111101101110100000010101000101001001110101001101110101101101010001101001000010110010000101111111100001010000010001100010001101000100;
XPCT = 108'b001111100101000001000110001001101000110011111010101110000000010000000110011000000000100000111110010001110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30600

pattern = 153; // 30600
ALLPIS = 207'b010000011010000011100011101011000110101110011010011100010110001000000100110100000110010011100010101000101110000110000011111011010011111010000001011111100010100110110010101111000010010010110100110011101001010;
XPCT = 108'b001101110001001001011010011011101001100011111001111110010000011110110100011001010110101101100111111111101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30800

pattern = 154; // 30800
ALLPIS = 207'b101001010100001011001101000000100110111001101110100011111101111101010111011100101100100000010111000011010010101011010100110101100110011010000001000111001011011010001000110111110011010011111000110001110111000;
XPCT = 108'b110110111001101001111100011001110111101011111110101111011001001000011110110111110000111111000001001010100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31000

pattern = 155; // 31000
ALLPIS = 207'b100001101010000001101010100000010001111111011110001111101110100110001101010101000001010101111011000110000110111100010000110111010001010110000001010000000110000000010001011110001111110000110001011010111111100;
XPCT = 108'b110011110111111000011000101110111111110011101111111111000110110111011111110000011001100000111110010010110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31200

pattern = 156; // 31200
ALLPIS = 207'b110101101101100000111001100110001110000101101101110011010010010111101110011101100111100001111001110010101001001111001000111010101000010010110110010111100111100001111101000010110101110101011100001100010011110;
XPCT = 108'b110000011010111010101110000100010011111111011111111111001111001111011111101111001000111010100111110110001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31400

pattern = 157; // 31400
ALLPIS = 207'b101001011100001001010100111000111011001010101111001101000000001111101011011110101011100110110111101100000101101010001010011011110111001101010101010011000011111011010000010001100011111101000001111101010101001;
XPCT = 108'b110010001001111110100000111101010101100101111111111111010110101000011111010011111110101010111111000101011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31600

pattern = 158; // 31600
ALLPIS = 207'b000011100010011110111011101101100101001101101110100011100000100010001111010011000001101000011011011000011000110001010100001110010000110111011110000000101100100100011101100111000111001100110001101100000101001;
XPCT = 108'b000100110011100110011000110100000101010111111010001010011001000011001110110100101001111111100001111110110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31800

pattern = 159; // 31800
ALLPIS = 207'b000100011110000100100010001101110110000101101000001100011001101110110010000001110010100010101011011110101111011111101001010001010101010100010101100001111110100101100001110000111000100110011110101111001110001;
XPCT = 108'b000110001100010011001111010111001110111101111001110100011111010010001111100101101010110110100000001100001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32000

pattern = 160; // 32000
ALLPIS = 207'b010101110011001110111010110010110011101010110010100111010010111010101111111011101100011000101000011101011100000000111011100110001111111001111101010001101011101101000100111101110111111011101010010011011100100;
XPCT = 108'b000111101011111101110101001011011100101011111011111110001111100001011111011111101000110110111000110000100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32200

pattern = 161; // 32200
ALLPIS = 207'b001001100101011101000110000110001000011100100110111111010110011010100011100001001110001111111010101000000010111000010100100111010111100100010101001001001111001100000001110011001101110101000111100000111000110;
XPCT = 108'b000110010110111010100011110000111000110001111011111110001111010001011111010100111001111001000001101001010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32400

pattern = 162; // 32400
ALLPIS = 207'b101000011001111110110101001001101111011011100011100101100110110001100011001101000000011011001011010100101111110111100111000011110000010100111110010010100111101111001011101001111100000011110101100000110111100;
XPCT = 108'b111101001110000001111010110000110111111001001110101111101111100000101111000101100100111111111111100110110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32600

pattern = 163; // 32600
ALLPIS = 207'b100010101110111111001010001001010101110011100111001100100111010001001110110101101011100101110010010011001101010001000000010001010011001011101001011001100001100001001010101011001001000001111100110000111011111;
XPCT = 108'b111101010100100000111110011000111011000011111100001011000000011011001110111001000110101111011001101000111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32800

pattern = 164; // 32800
ALLPIS = 207'b010101110110010111110101101100101000110111000100100011110100011000101101010100111101100010011101010010010101001100101010110000011010011110100101110010011011110001010001101101101001100010010110010011010100010;
XPCT = 108'b000101101100110001001011001011010100110010111011111110010000011001011110010001001110100010011000111010010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33000

pattern = 165; // 33000
ALLPIS = 207'b011110010010111100000111011100110000100000110101001011111111111011111000010111000110110111000100100100010101110100100101000110100100000010010100010111001001111110011011101001111000111110010011001010111010010;
XPCT = 108'b001101001100011111001001100110111010011011111011011010000000100000001110101000100100100001111110000000000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33200

pattern = 166; // 33200
ALLPIS = 207'b000110100100000011101111010011000001111010010010110111110100010001000000011011101001111000100010101100110011010111110010001011010110010010000110111101100101001001000000110001000001111110011010100010010011100;
XPCT = 108'b000110000000111111001101010010010011000011111011011010001111011001001111101111111000111111100001001110100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33400

pattern = 167; // 33400
ALLPIS = 207'b111111000100010000111101010011100011010110010110101000101000111011001000101000110010110001010010001111100001000111000101101001000010001000010000101100011110010111011011000110101000000001001001100111100100100;
XPCT = 108'b111000111100000000100100110011100100010111111101011011000000001100111110111000011111100000111110100000010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33600

pattern = 168; // 33600
ALLPIS = 207'b010110100110100001010100101111000110000110011100011001100111010111000110110000111010110110110100010110010011111110000111010101010101000100111100110111100111001010110100110011101101111100011111111010110001000;
XPCT = 108'b000110011110111110001111111110110001000011111011011010001111011001111111101111101000111111000000110001010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33800

pattern = 169; // 33800
ALLPIS = 207'b100000101100101111101111010000101111011000000000010101010000010000000100101011000111011100111111101101001000111110001010111010011100001101001111000110101001000100110110000101010010100110010111011101110110101;
XPCT = 108'b111000100001010011001011101101110110101111110111111111111111101111001111111101001101110110100001011111111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34000

pattern = 170; // 34000
ALLPIS = 207'b101100110110000000001011101001010010110110010111110100111111101000101100101101001110101100100010100111111110110111110100100010000110111000101101110101100000011110111111010101001000000111010011101110011010111;
XPCT = 108'b111010100100000011101001110110011010110111101100101111110000001100011110101001001011101000111001100010101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34200

pattern = 171; // 34200
ALLPIS = 207'b100000110110111101110100000010100101101100110100001100000000011001100001111000011110100010110111010101011111110110101010101110001111010001000011110000000011101101110000110001000001000010110100110001000001100;
XPCT = 108'b110110000000100001011010011001000001100001101101111111011111101111001111010100101010111111000001011111100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34400

pattern = 172; // 34400
ALLPIS = 207'b110110011001011010001110010010101000101100010111010010100001010011011011000010010100110010110000010011010010000101100100011000011001010101100010000001011100110000010000010100110101110010110011001101010000101;
XPCT = 108'b110010101010111001011001100101010000001111111101011011001111100000001111110100111011111100011110000000001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34600

pattern = 173; // 34600
ALLPIS = 207'b011001011001011101100110010111001001010001110000010001101101100011111111010100110100100110011101101101011011000000000001010111101111100000000000101101010111101001110011100110011000100101111100011000001000010;
XPCT = 108'b001100110100010010111110001100001000111010111011111110010110100101011111110000101100101010011111101000110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34800

pattern = 174; // 34800
ALLPIS = 207'b101011110011110101101111100110101100101110000111011100111001111101011100000011111001000010100001100101101000111110110001011110010110110111001000100010110001111101111100101001011101010001111000011010101101000;
XPCT = 108'b110101000110101000111100001110101101001011111100001011011111010111111111010111010011111100011111101011000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35000

pattern = 175; // 35000
ALLPIS = 207'b011011011100111111000111110100000110010000011101001111001111100101110110000101000011001111010111101110000101100100001010111010110110101101001110111011001010110100010111001111101100101100110111010011010000010;
XPCT = 108'b001001111110010110011011101011010000010011111011011010010000100011111110010000001001100111000000000101100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35200

pattern = 176; // 35200
ALLPIS = 207'b110100111000101011100111111110111001011000110111000010101100111101100011010000000110000000110001000111010001000010110011010001010000000100100100010101000010111110001000000001010111100101011010101001000010000;
XPCT = 108'b110000000011110010101101010101000010101011111101111111011111100000001011010110111111110101100001010110000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35400

pattern = 177; // 35400
ALLPIS = 207'b011001001000000100011001011011001011011100011100101000011000011011001111111011001111000010001010100011001001100011000001110110100001110101111101000100010011011101110011100010110000000100000111111111100011101;
XPCT = 108'b001100011000000010000011111111100011111110111001111110001111010111100111100111100110110100100001100011101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35600

pattern = 178; // 35600
ALLPIS = 207'b000111001000011110100100110101110000001011010001111001011101100000110000000100111101110100010110101111001110001001110010100000111101001110010000011111100011110011000111000101000011110110100011010010111000010;
XPCT = 108'b001000100001111011010001101010111000010001111011010000010110000101001111001000010110101000011110010000011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35800

pattern = 179; // 35800
ALLPIS = 207'b100011100100001111010010011010111000000101101000111100101110110000011000000010011110111010001011010111100111000100111001010000011110100111001000001111110001111001100011100010100001111011010001101001011100001;
XPCT = 108'b111100011000111101101000110101011100010001111101011011111001011000011110100101011011110010100000101110110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36000

pattern = 180; // 36000
ALLPIS = 207'b000010111000101000111111101011100101101011011001100100011000100000101010010010010101000100001101111101101011101000010101001000110110110000010101100001111110101010010110100111101100101111011001111001100110101;
XPCT = 108'b001100111110010111101100111101100110000010111001011010001111000110100101010110011110110010100000001001001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36200

      $display("// %t : Simulation of %0d patterns completed with %0d errors\n", $time, pattern+1, nofails);
      if (verbose >=2) $finish(2);
      /* else */ $finish(0);
   end
endmodule
