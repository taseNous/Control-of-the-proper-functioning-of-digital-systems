// Verilog pattern output written by  TetraMAX (TM)  B-2008.09-SP2-i081128_181834 
// Date: Wed Jul  6 12:10:26 2011
// Module tested: c7552

//     Uncollapsed Stuck Fault Summary Report
// -----------------------------------------------
// fault class                     code   #faults
// ------------------------------  ----  ---------
// Detected                         DT       6593
// Possibly detected                PT          0
// Undetectable                     UD          0
// ATPG untestable                  AU          0
// Not detected                     ND        295
// -----------------------------------------------
// total faults                              6888
// test coverage                            95.72%
// -----------------------------------------------
// 
//            Pattern Summary Report
// -----------------------------------------------
// #internal patterns                         175
//     #basic_scan patterns                   175
// -----------------------------------------------
// 
// There are no rule fails
// There are no clocks
// There are no constraint ports
// There are no equivalent pins
// There are no net connections

`timescale 1 ns / 1 ns

//
// --- NOTE: Remove the comment to define 'tmax_iddq' to activate processing of IDDQ events
//     Or use '+define+tmax_iddq' on the verilog compile line
//
//`define tmax_iddq

module AAA_tmax_testbench_1_16 ;
   parameter NAMELENGTH = 200; // max length of names reported in fails
   integer nofails, bit, pattern, lastpattern;
   integer error_banner; // flag for tracking displayed error banner
   integer loads;        // number of load_unloads for current pattern
   integer patm1;        // pattern - 1
   integer patp1;        // pattern + lastpattern
   integer prev_pat;     // previous pattern number
   integer report_interval; // report pattern progress every Nth pattern
   integer verbose;      // message verbosity level
   parameter NINPUTS = 207, NOUTPUTS = 108;
   wire [0:NOUTPUTS-1] PO; reg [0:NOUTPUTS-1] ALLPOS, XPCT, MASK;
   reg [0:NINPUTS-1] PI, ALLPIS;
   reg [0:8*(NAMELENGTH-1)] POnames [0:NOUTPUTS-1];
   event IDDQ;

   wire N1;
   wire N5;
   wire N9;
   wire N12;
   wire N15;
   wire N18;
   wire N23;
   wire N26;
   wire N29;
   wire N32;
   wire N35;
   wire N38;
   wire N41;
   wire N44;
   wire N47;
   wire N50;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N69;
   wire N70;
   wire N73;
   wire N74;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N82;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N94;
   wire N97;
   wire N100;
   wire N103;
   wire N106;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N118;
   wire N121;
   wire N124;
   wire N127;
   wire N130;
   wire N133;
   wire N134;
   wire N135;
   wire N138;
   wire N141;
   wire N144;
   wire N147;
   wire N150;
   wire N151;
   wire N152;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N178;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire N185;
   wire N186;
   wire N187;
   wire N188;
   wire N189;
   wire N190;
   wire N191;
   wire N192;
   wire N193;
   wire N194;
   wire N195;
   wire N196;
   wire N197;
   wire N198;
   wire N199;
   wire N200;
   wire N201;
   wire N202;
   wire N203;
   wire N204;
   wire N205;
   wire N206;
   wire N207;
   wire N208;
   wire N209;
   wire N210;
   wire N211;
   wire N212;
   wire N213;
   wire N214;
   wire N215;
   wire N216;
   wire N217;
   wire N218;
   wire N219;
   wire N220;
   wire N221;
   wire N222;
   wire N223;
   wire N224;
   wire N225;
   wire N226;
   wire N227;
   wire N228;
   wire N229;
   wire N230;
   wire N231;
   wire N232;
   wire N233;
   wire N234;
   wire N235;
   wire N236;
   wire N237;
   wire N238;
   wire N239;
   wire N240;
   wire N242;
   wire N245;
   wire N248;
   wire N251;
   wire N254;
   wire N257;
   wire N260;
   wire N263;
   wire N267;
   wire N271;
   wire N274;
   wire N277;
   wire N280;
   wire N283;
   wire N286;
   wire N289;
   wire N293;
   wire N296;
   wire N299;
   wire N303;
   wire N307;
   wire N310;
   wire N313;
   wire N316;
   wire N319;
   wire N322;
   wire N325;
   wire N328;
   wire N331;
   wire N334;
   wire N337;
   wire N340;
   wire N343;
   wire N346;
   wire N349;
   wire N352;
   wire N355;
   wire N358;
   wire N361;
   wire N364;
   wire N367;
   wire N382;
   wire N241_I;
   wire N387;
   wire N388;
   wire N478;
   wire N482;
   wire N484;
   wire N486;
   wire N489;
   wire N492;
   wire N501;
   wire N505;
   wire N507;
   wire N509;
   wire N511;
   wire N513;
   wire N515;
   wire N517;
   wire N519;
   wire N535;
   wire N537;
   wire N539;
   wire N541;
   wire N543;
   wire N545;
   wire N547;
   wire N549;
   wire N551;
   wire N553;
   wire N556;
   wire N559;
   wire N561;
   wire N563;
   wire N565;
   wire N567;
   wire N569;
   wire N571;
   wire N573;
   wire N582;
   wire N643;
   wire N707;
   wire N813;
   wire N881;
   wire N882;
   wire N883;
   wire N884;
   wire N885;
   wire N889;
   wire N945;
   wire N1110;
   wire N1111;
   wire N1112;
   wire N1113;
   wire N1114;
   wire N1489;
   wire N1490;
   wire N1781;
   wire N10025;
   wire N10101;
   wire N10102;
   wire N10103;
   wire N10104;
   wire N10109;
   wire N10110;
   wire N10111;
   wire N10112;
   wire N10350;
   wire N10351;
   wire N10352;
   wire N10353;
   wire N10574;
   wire N10575;
   wire N10576;
   wire N10628;
   wire N10632;
   wire N10641;
   wire N10704;
   wire N10706;
   wire N10711;
   wire N10712;
   wire N10713;
   wire N10714;
   wire N10715;
   wire N10716;
   wire N10717;
   wire N10718;
   wire N10729;
   wire N10759;
   wire N10760;
   wire N10761;
   wire N10762;
   wire N10763;
   wire N10827;
   wire N10837;
   wire N10838;
   wire N10839;
   wire N10840;
   wire N10868;
   wire N10869;
   wire N10870;
   wire N10871;
   wire N10905;
   wire N10906;
   wire N10907;
   wire N10908;
   wire N11333;
   wire N11334;
   wire N11340;
   wire N11342;
   wire N241_O;

   // map PI[] vector to DUT inputs and bidis
   assign N1 = PI[0];
   assign N5 = PI[1];
   assign N9 = PI[2];
   assign N12 = PI[3];
   assign N15 = PI[4];
   assign N18 = PI[5];
   assign N23 = PI[6];
   assign N26 = PI[7];
   assign N29 = PI[8];
   assign N32 = PI[9];
   assign N35 = PI[10];
   assign N38 = PI[11];
   assign N41 = PI[12];
   assign N44 = PI[13];
   assign N47 = PI[14];
   assign N50 = PI[15];
   assign N53 = PI[16];
   assign N54 = PI[17];
   assign N55 = PI[18];
   assign N56 = PI[19];
   assign N57 = PI[20];
   assign N58 = PI[21];
   assign N59 = PI[22];
   assign N60 = PI[23];
   assign N61 = PI[24];
   assign N62 = PI[25];
   assign N63 = PI[26];
   assign N64 = PI[27];
   assign N65 = PI[28];
   assign N66 = PI[29];
   assign N69 = PI[30];
   assign N70 = PI[31];
   assign N73 = PI[32];
   assign N74 = PI[33];
   assign N75 = PI[34];
   assign N76 = PI[35];
   assign N77 = PI[36];
   assign N78 = PI[37];
   assign N79 = PI[38];
   assign N80 = PI[39];
   assign N81 = PI[40];
   assign N82 = PI[41];
   assign N83 = PI[42];
   assign N84 = PI[43];
   assign N85 = PI[44];
   assign N86 = PI[45];
   assign N87 = PI[46];
   assign N88 = PI[47];
   assign N89 = PI[48];
   assign N94 = PI[49];
   assign N97 = PI[50];
   assign N100 = PI[51];
   assign N103 = PI[52];
   assign N106 = PI[53];
   assign N109 = PI[54];
   assign N110 = PI[55];
   assign N111 = PI[56];
   assign N112 = PI[57];
   assign N113 = PI[58];
   assign N114 = PI[59];
   assign N115 = PI[60];
   assign N118 = PI[61];
   assign N121 = PI[62];
   assign N124 = PI[63];
   assign N127 = PI[64];
   assign N130 = PI[65];
   assign N133 = PI[66];
   assign N134 = PI[67];
   assign N135 = PI[68];
   assign N138 = PI[69];
   assign N141 = PI[70];
   assign N144 = PI[71];
   assign N147 = PI[72];
   assign N150 = PI[73];
   assign N151 = PI[74];
   assign N152 = PI[75];
   assign N153 = PI[76];
   assign N154 = PI[77];
   assign N155 = PI[78];
   assign N156 = PI[79];
   assign N157 = PI[80];
   assign N158 = PI[81];
   assign N159 = PI[82];
   assign N160 = PI[83];
   assign N161 = PI[84];
   assign N162 = PI[85];
   assign N163 = PI[86];
   assign N164 = PI[87];
   assign N165 = PI[88];
   assign N166 = PI[89];
   assign N167 = PI[90];
   assign N168 = PI[91];
   assign N169 = PI[92];
   assign N170 = PI[93];
   assign N171 = PI[94];
   assign N172 = PI[95];
   assign N173 = PI[96];
   assign N174 = PI[97];
   assign N175 = PI[98];
   assign N176 = PI[99];
   assign N177 = PI[100];
   assign N178 = PI[101];
   assign N179 = PI[102];
   assign N180 = PI[103];
   assign N181 = PI[104];
   assign N182 = PI[105];
   assign N183 = PI[106];
   assign N184 = PI[107];
   assign N185 = PI[108];
   assign N186 = PI[109];
   assign N187 = PI[110];
   assign N188 = PI[111];
   assign N189 = PI[112];
   assign N190 = PI[113];
   assign N191 = PI[114];
   assign N192 = PI[115];
   assign N193 = PI[116];
   assign N194 = PI[117];
   assign N195 = PI[118];
   assign N196 = PI[119];
   assign N197 = PI[120];
   assign N198 = PI[121];
   assign N199 = PI[122];
   assign N200 = PI[123];
   assign N201 = PI[124];
   assign N202 = PI[125];
   assign N203 = PI[126];
   assign N204 = PI[127];
   assign N205 = PI[128];
   assign N206 = PI[129];
   assign N207 = PI[130];
   assign N208 = PI[131];
   assign N209 = PI[132];
   assign N210 = PI[133];
   assign N211 = PI[134];
   assign N212 = PI[135];
   assign N213 = PI[136];
   assign N214 = PI[137];
   assign N215 = PI[138];
   assign N216 = PI[139];
   assign N217 = PI[140];
   assign N218 = PI[141];
   assign N219 = PI[142];
   assign N220 = PI[143];
   assign N221 = PI[144];
   assign N222 = PI[145];
   assign N223 = PI[146];
   assign N224 = PI[147];
   assign N225 = PI[148];
   assign N226 = PI[149];
   assign N227 = PI[150];
   assign N228 = PI[151];
   assign N229 = PI[152];
   assign N230 = PI[153];
   assign N231 = PI[154];
   assign N232 = PI[155];
   assign N233 = PI[156];
   assign N234 = PI[157];
   assign N235 = PI[158];
   assign N236 = PI[159];
   assign N237 = PI[160];
   assign N238 = PI[161];
   assign N239 = PI[162];
   assign N240 = PI[163];
   assign N242 = PI[164];
   assign N245 = PI[165];
   assign N248 = PI[166];
   assign N251 = PI[167];
   assign N254 = PI[168];
   assign N257 = PI[169];
   assign N260 = PI[170];
   assign N263 = PI[171];
   assign N267 = PI[172];
   assign N271 = PI[173];
   assign N274 = PI[174];
   assign N277 = PI[175];
   assign N280 = PI[176];
   assign N283 = PI[177];
   assign N286 = PI[178];
   assign N289 = PI[179];
   assign N293 = PI[180];
   assign N296 = PI[181];
   assign N299 = PI[182];
   assign N303 = PI[183];
   assign N307 = PI[184];
   assign N310 = PI[185];
   assign N313 = PI[186];
   assign N316 = PI[187];
   assign N319 = PI[188];
   assign N322 = PI[189];
   assign N325 = PI[190];
   assign N328 = PI[191];
   assign N331 = PI[192];
   assign N334 = PI[193];
   assign N337 = PI[194];
   assign N340 = PI[195];
   assign N343 = PI[196];
   assign N346 = PI[197];
   assign N349 = PI[198];
   assign N352 = PI[199];
   assign N355 = PI[200];
   assign N358 = PI[201];
   assign N361 = PI[202];
   assign N364 = PI[203];
   assign N367 = PI[204];
   assign N382 = PI[205];
   assign N241_I = PI[206];

   // map DUT outputs and bidis to PO[] vector
   assign
      PO[0] = N387 ,
      PO[1] = N388 ,
      PO[2] = N478 ,
      PO[3] = N482 ,
      PO[4] = N484 ,
      PO[5] = N486 ,
      PO[6] = N489 ,
      PO[7] = N492 ,
      PO[8] = N501 ,
      PO[9] = N505 ,
      PO[10] = N507 ,
      PO[11] = N509 ,
      PO[12] = N511 ,
      PO[13] = N513 ,
      PO[14] = N515 ,
      PO[15] = N517 ,
      PO[16] = N519 ,
      PO[17] = N535 ,
      PO[18] = N537 ,
      PO[19] = N539 ,
      PO[20] = N541 ,
      PO[21] = N543 ,
      PO[22] = N545 ,
      PO[23] = N547 ,
      PO[24] = N549 ,
      PO[25] = N551 ,
      PO[26] = N553 ,
      PO[27] = N556 ,
      PO[28] = N559 ,
      PO[29] = N561 ,
      PO[30] = N563 ,
      PO[31] = N565 ;
   assign
      PO[32] = N567 ,
      PO[33] = N569 ,
      PO[34] = N571 ,
      PO[35] = N573 ,
      PO[36] = N582 ,
      PO[37] = N643 ,
      PO[38] = N707 ,
      PO[39] = N813 ,
      PO[40] = N881 ,
      PO[41] = N882 ,
      PO[42] = N883 ,
      PO[43] = N884 ,
      PO[44] = N885 ,
      PO[45] = N889 ,
      PO[46] = N945 ,
      PO[47] = N1110 ,
      PO[48] = N1111 ,
      PO[49] = N1112 ,
      PO[50] = N1113 ,
      PO[51] = N1114 ,
      PO[52] = N1489 ,
      PO[53] = N1490 ,
      PO[54] = N1781 ,
      PO[55] = N10025 ,
      PO[56] = N10101 ,
      PO[57] = N10102 ,
      PO[58] = N10103 ,
      PO[59] = N10104 ,
      PO[60] = N10109 ,
      PO[61] = N10110 ,
      PO[62] = N10111 ,
      PO[63] = N10112 ;
   assign
      PO[64] = N10350 ,
      PO[65] = N10351 ,
      PO[66] = N10352 ,
      PO[67] = N10353 ,
      PO[68] = N10574 ,
      PO[69] = N10575 ,
      PO[70] = N10576 ,
      PO[71] = N10628 ,
      PO[72] = N10632 ,
      PO[73] = N10641 ,
      PO[74] = N10704 ,
      PO[75] = N10706 ,
      PO[76] = N10711 ,
      PO[77] = N10712 ,
      PO[78] = N10713 ,
      PO[79] = N10714 ,
      PO[80] = N10715 ,
      PO[81] = N10716 ,
      PO[82] = N10717 ,
      PO[83] = N10718 ,
      PO[84] = N10729 ,
      PO[85] = N10759 ,
      PO[86] = N10760 ,
      PO[87] = N10761 ,
      PO[88] = N10762 ,
      PO[89] = N10763 ,
      PO[90] = N10827 ,
      PO[91] = N10837 ,
      PO[92] = N10838 ,
      PO[93] = N10839 ,
      PO[94] = N10840 ,
      PO[95] = N10868 ;
   assign
      PO[96] = N10869 ,
      PO[97] = N10870 ,
      PO[98] = N10871 ,
      PO[99] = N10905 ,
      PO[100] = N10906 ,
      PO[101] = N10907 ,
      PO[102] = N10908 ,
      PO[103] = N11333 ,
      PO[104] = N11334 ,
      PO[105] = N11340 ,
      PO[106] = N11342 ,
      PO[107] = N241_O ;

   // instantiate the design into the testbench
   c7552 dut (
      .N1(N1),
      .N5(N5),
      .N9(N9),
      .N12(N12),
      .N15(N15),
      .N18(N18),
      .N23(N23),
      .N26(N26),
      .N29(N29),
      .N32(N32),
      .N35(N35),
      .N38(N38),
      .N41(N41),
      .N44(N44),
      .N47(N47),
      .N50(N50),
      .N53(N53),
      .N54(N54),
      .N55(N55),
      .N56(N56),
      .N57(N57),
      .N58(N58),
      .N59(N59),
      .N60(N60),
      .N61(N61),
      .N62(N62),
      .N63(N63),
      .N64(N64),
      .N65(N65),
      .N66(N66),
      .N69(N69),
      .N70(N70),
      .N73(N73),
      .N74(N74),
      .N75(N75),
      .N76(N76),
      .N77(N77),
      .N78(N78),
      .N79(N79),
      .N80(N80),
      .N81(N81),
      .N82(N82),
      .N83(N83),
      .N84(N84),
      .N85(N85),
      .N86(N86),
      .N87(N87),
      .N88(N88),
      .N89(N89),
      .N94(N94),
      .N97(N97),
      .N100(N100),
      .N103(N103),
      .N106(N106),
      .N109(N109),
      .N110(N110),
      .N111(N111),
      .N112(N112),
      .N113(N113),
      .N114(N114),
      .N115(N115),
      .N118(N118),
      .N121(N121),
      .N124(N124),
      .N127(N127),
      .N130(N130),
      .N133(N133),
      .N134(N134),
      .N135(N135),
      .N138(N138),
      .N141(N141),
      .N144(N144),
      .N147(N147),
      .N150(N150),
      .N151(N151),
      .N152(N152),
      .N153(N153),
      .N154(N154),
      .N155(N155),
      .N156(N156),
      .N157(N157),
      .N158(N158),
      .N159(N159),
      .N160(N160),
      .N161(N161),
      .N162(N162),
      .N163(N163),
      .N164(N164),
      .N165(N165),
      .N166(N166),
      .N167(N167),
      .N168(N168),
      .N169(N169),
      .N170(N170),
      .N171(N171),
      .N172(N172),
      .N173(N173),
      .N174(N174),
      .N175(N175),
      .N176(N176),
      .N177(N177),
      .N178(N178),
      .N179(N179),
      .N180(N180),
      .N181(N181),
      .N182(N182),
      .N183(N183),
      .N184(N184),
      .N185(N185),
      .N186(N186),
      .N187(N187),
      .N188(N188),
      .N189(N189),
      .N190(N190),
      .N191(N191),
      .N192(N192),
      .N193(N193),
      .N194(N194),
      .N195(N195),
      .N196(N196),
      .N197(N197),
      .N198(N198),
      .N199(N199),
      .N200(N200),
      .N201(N201),
      .N202(N202),
      .N203(N203),
      .N204(N204),
      .N205(N205),
      .N206(N206),
      .N207(N207),
      .N208(N208),
      .N209(N209),
      .N210(N210),
      .N211(N211),
      .N212(N212),
      .N213(N213),
      .N214(N214),
      .N215(N215),
      .N216(N216),
      .N217(N217),
      .N218(N218),
      .N219(N219),
      .N220(N220),
      .N221(N221),
      .N222(N222),
      .N223(N223),
      .N224(N224),
      .N225(N225),
      .N226(N226),
      .N227(N227),
      .N228(N228),
      .N229(N229),
      .N230(N230),
      .N231(N231),
      .N232(N232),
      .N233(N233),
      .N234(N234),
      .N235(N235),
      .N236(N236),
      .N237(N237),
      .N238(N238),
      .N239(N239),
      .N240(N240),
      .N242(N242),
      .N245(N245),
      .N248(N248),
      .N251(N251),
      .N254(N254),
      .N257(N257),
      .N260(N260),
      .N263(N263),
      .N267(N267),
      .N271(N271),
      .N274(N274),
      .N277(N277),
      .N280(N280),
      .N283(N283),
      .N286(N286),
      .N289(N289),
      .N293(N293),
      .N296(N296),
      .N299(N299),
      .N303(N303),
      .N307(N307),
      .N310(N310),
      .N313(N313),
      .N316(N316),
      .N319(N319),
      .N322(N322),
      .N325(N325),
      .N328(N328),
      .N331(N331),
      .N334(N334),
      .N337(N337),
      .N340(N340),
      .N343(N343),
      .N346(N346),
      .N349(N349),
      .N352(N352),
      .N355(N355),
      .N358(N358),
      .N361(N361),
      .N364(N364),
      .N367(N367),
      .N382(N382),
      .N241_I(N241_I),
      .N387(N387),
      .N388(N388),
      .N478(N478),
      .N482(N482),
      .N484(N484),
      .N486(N486),
      .N489(N489),
      .N492(N492),
      .N501(N501),
      .N505(N505),
      .N507(N507),
      .N509(N509),
      .N511(N511),
      .N513(N513),
      .N515(N515),
      .N517(N517),
      .N519(N519),
      .N535(N535),
      .N537(N537),
      .N539(N539),
      .N541(N541),
      .N543(N543),
      .N545(N545),
      .N547(N547),
      .N549(N549),
      .N551(N551),
      .N553(N553),
      .N556(N556),
      .N559(N559),
      .N561(N561),
      .N563(N563),
      .N565(N565),
      .N567(N567),
      .N569(N569),
      .N571(N571),
      .N573(N573),
      .N582(N582),
      .N643(N643),
      .N707(N707),
      .N813(N813),
      .N881(N881),
      .N882(N882),
      .N883(N883),
      .N884(N884),
      .N885(N885),
      .N889(N889),
      .N945(N945),
      .N1110(N1110),
      .N1111(N1111),
      .N1112(N1112),
      .N1113(N1113),
      .N1114(N1114),
      .N1489(N1489),
      .N1490(N1490),
      .N1781(N1781),
      .N10025(N10025),
      .N10101(N10101),
      .N10102(N10102),
      .N10103(N10103),
      .N10104(N10104),
      .N10109(N10109),
      .N10110(N10110),
      .N10111(N10111),
      .N10112(N10112),
      .N10350(N10350),
      .N10351(N10351),
      .N10352(N10352),
      .N10353(N10353),
      .N10574(N10574),
      .N10575(N10575),
      .N10576(N10576),
      .N10628(N10628),
      .N10632(N10632),
      .N10641(N10641),
      .N10704(N10704),
      .N10706(N10706),
      .N10711(N10711),
      .N10712(N10712),
      .N10713(N10713),
      .N10714(N10714),
      .N10715(N10715),
      .N10716(N10716),
      .N10717(N10717),
      .N10718(N10718),
      .N10729(N10729),
      .N10759(N10759),
      .N10760(N10760),
      .N10761(N10761),
      .N10762(N10762),
      .N10763(N10763),
      .N10827(N10827),
      .N10837(N10837),
      .N10838(N10838),
      .N10839(N10839),
      .N10840(N10840),
      .N10868(N10868),
      .N10869(N10869),
      .N10870(N10870),
      .N10871(N10871),
      .N10905(N10905),
      .N10906(N10906),
      .N10907(N10907),
      .N10908(N10908),
      .N11333(N11333),
      .N11334(N11334),
      .N11340(N11340),
      .N11342(N11342),
      .N241_O(N241_O)   );


   integer errshown;
   event measurePO;
   always @ measurePO begin
      if (((XPCT&MASK) !== (ALLPOS&MASK)) || (XPCT !== (~(~XPCT)))) begin
         errshown = 0;
         for (bit = 0; bit < NOUTPUTS; bit=bit + 1) begin
            if (MASK[bit]==1'b1) begin
               if (XPCT[bit] !== ALLPOS[bit]) begin
                  if (errshown==0) $display("\n// *** ERROR during capture pattern %0d, T=%t", pattern, $time);
                  $display("  %0d %0s (exp=%b, got=%b)", pattern, POnames[bit], XPCT[bit], ALLPOS[bit]);
                  nofails = nofails + 1; errshown = 1;
               end
            end
         end
      end
   end

   event forcePI_default_WFT;
   always @ forcePI_default_WFT begin
      PI = ALLPIS;
   end
   event measurePO_default_WFT;
   always @ measurePO_default_WFT begin
      #40;
      ALLPOS = PO;
      #0; #0 -> measurePO;
      `ifdef tmax_iddq
         #0; ->IDDQ;
      `endif
   end

   always @ IDDQ begin
   `ifdef tmax_iddq
      $ssi_iddq("strobe_try");
      $ssi_iddq("status drivers leaky AAA_tmax_testbench_1_16.leaky");
   `endif
   end

   event capture;
   always @ capture begin
      ->forcePI_default_WFT;
      #100; ->measurePO_default_WFT;
   end


   initial begin

      //
      // --- establish a default time format for %t
      //
      $timeformat(-9,2," ns",18);

      //
      // --- default verbosity to 2 but also allow user override by
      //     using '+define+tmax_msg=N' on verilog compile line.
      //
      `ifdef tmax_msg
         verbose = `tmax_msg ;
      `else
         verbose = 2 ;
      `endif

      //
      // --- default pattern reporting interval to 5 but also allow user
      //     override by using '+define+tmax_rpt=N' on verilog compile line.
      //
      `ifdef tmax_rpt
         report_interval = `tmax_rpt ;
      `else
         report_interval = 5 ;
      `endif

      //
      // --- support generating Extened VCD output by using
      //     '+define+tmax_vcde' on verilog compile line.
      //
      `ifdef tmax_vcde
         // extended VCD, see IEEE Verilog P1364.1-1999 Draft 2
         if (verbose >= 2) $display("// %t : opening Extended VCD output file", $time);
         $dumpports( dut, "sim_vcde.out");
      `endif

      //
      // --- IDDQ PLI initialization
      //     User may activite by using '+define+tmax_iddq' on verilog compile line.
      //     Or by defining `tmax_iddq in this file.
      //
      `ifdef tmax_iddq
         if (verbose >= 3) $display("// %t : Initializing IDDQ PLI", $time);
         $ssi_iddq("dut AAA_tmax_testbench_1_16.dut");
         $ssi_iddq("verb on");
         $ssi_iddq("cycle 0");
         //
         // --- User may select one of the following two methods for fault seeding:
         //     #1 faults seeded by PLI (default)
         //     #2 faults supplied in a file
         //     Comment out the unused lines as needed (precede with '//').
         //     Replace the 'FAULTLIST_FILE' string with the actual file pathname.
         //
         $ssi_iddq("seed SA AAA_tmax_testbench_1_16.dut");   // no file, faults seeded by PLI
         //
         // $ssi_iddq("scope AAA_tmax_testbench_1_16.dut");   // set scope for faults from a file
         // $ssi_iddq("read_tmax FAULTLIST_FILE"); // read faults from a file
         //
      `endif

      POnames[0] = "N387";
      POnames[1] = "N388";
      POnames[2] = "N478";
      POnames[3] = "N482";
      POnames[4] = "N484";
      POnames[5] = "N486";
      POnames[6] = "N489";
      POnames[7] = "N492";
      POnames[8] = "N501";
      POnames[9] = "N505";
      POnames[10] = "N507";
      POnames[11] = "N509";
      POnames[12] = "N511";
      POnames[13] = "N513";
      POnames[14] = "N515";
      POnames[15] = "N517";
      POnames[16] = "N519";
      POnames[17] = "N535";
      POnames[18] = "N537";
      POnames[19] = "N539";
      POnames[20] = "N541";
      POnames[21] = "N543";
      POnames[22] = "N545";
      POnames[23] = "N547";
      POnames[24] = "N549";
      POnames[25] = "N551";
      POnames[26] = "N553";
      POnames[27] = "N556";
      POnames[28] = "N559";
      POnames[29] = "N561";
      POnames[30] = "N563";
      POnames[31] = "N565";
      POnames[32] = "N567";
      POnames[33] = "N569";
      POnames[34] = "N571";
      POnames[35] = "N573";
      POnames[36] = "N582";
      POnames[37] = "N643";
      POnames[38] = "N707";
      POnames[39] = "N813";
      POnames[40] = "N881";
      POnames[41] = "N882";
      POnames[42] = "N883";
      POnames[43] = "N884";
      POnames[44] = "N885";
      POnames[45] = "N889";
      POnames[46] = "N945";
      POnames[47] = "N1110";
      POnames[48] = "N1111";
      POnames[49] = "N1112";
      POnames[50] = "N1113";
      POnames[51] = "N1114";
      POnames[52] = "N1489";
      POnames[53] = "N1490";
      POnames[54] = "N1781";
      POnames[55] = "N10025";
      POnames[56] = "N10101";
      POnames[57] = "N10102";
      POnames[58] = "N10103";
      POnames[59] = "N10104";
      POnames[60] = "N10109";
      POnames[61] = "N10110";
      POnames[62] = "N10111";
      POnames[63] = "N10112";
      POnames[64] = "N10350";
      POnames[65] = "N10351";
      POnames[66] = "N10352";
      POnames[67] = "N10353";
      POnames[68] = "N10574";
      POnames[69] = "N10575";
      POnames[70] = "N10576";
      POnames[71] = "N10628";
      POnames[72] = "N10632";
      POnames[73] = "N10641";
      POnames[74] = "N10704";
      POnames[75] = "N10706";
      POnames[76] = "N10711";
      POnames[77] = "N10712";
      POnames[78] = "N10713";
      POnames[79] = "N10714";
      POnames[80] = "N10715";
      POnames[81] = "N10716";
      POnames[82] = "N10717";
      POnames[83] = "N10718";
      POnames[84] = "N10729";
      POnames[85] = "N10759";
      POnames[86] = "N10760";
      POnames[87] = "N10761";
      POnames[88] = "N10762";
      POnames[89] = "N10763";
      POnames[90] = "N10827";
      POnames[91] = "N10837";
      POnames[92] = "N10838";
      POnames[93] = "N10839";
      POnames[94] = "N10840";
      POnames[95] = "N10868";
      POnames[96] = "N10869";
      POnames[97] = "N10870";
      POnames[98] = "N10871";
      POnames[99] = "N10905";
      POnames[100] = "N10906";
      POnames[101] = "N10907";
      POnames[102] = "N10908";
      POnames[103] = "N11333";
      POnames[104] = "N11334";
      POnames[105] = "N11340";
      POnames[106] = "N11342";
      POnames[107] = "N241_O";
      nofails = 0; pattern = -1; lastpattern = 0;
      prev_pat = -2; error_banner = -2;
      /*** No test setup procedure ***/


      /*** Non-scan test ***/

      if (verbose >= 1) $display("// %t : Begin patterns, first pattern = 0", $time);
pattern = 0; // 0
ALLPIS = 207'b111010100010111101011100111110000111010001001110101011100001100110110110011011000100110110011111100111100111111110101101011001010100011101010110011010000001111111110110100011000110100111111111101000011100011;
XPCT = 108'b111100010011010011111111110100011100000011100111011011010110110011101111011000111100100110111000000001011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 200

pattern = 1; // 200
ALLPIS = 207'b011101010001011110101110011111000011101000100111010101110000110011011011001101100010011011001111110011110011111111010110101100101010001110101011001101000000111111111011010001100011010011111111110100001110001;
XPCT = 108'b001010001001101001111111111000001110110111110011111110011111111100111111101101101001111101111001100010110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 400

pattern = 2; // 400
ALLPIS = 207'b010100001010010010001011110001100110100101011101000001011001111111011011111101110101111011111000011110011110000001000110001111000001011010000011111100100001100000001011001011110111001110000000010010011011011;
XPCT = 108'b001001011011100111000000001010011011111011111011111110010000000011110100101011110101100010011001011101110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 600

pattern = 3; // 600
ALLPIS = 207'b110000100111110100011001000110110100000011100000001011001101011001011011100101111110001011100011101000101000111110001110011110110100110000010111100100010001001111110011000110111101000000111111100001010001110;
XPCT = 108'b111000111110100000011111110001010001111011111111111111111111110110011111100100101101111111000001011111010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 800

pattern = 4; // 800
ALLPIS = 207'b100010110001000111010000011101011101010000111110101110000111001010011011101001111011110011101110010011110011100001101010010110001110000101011101101000001001011000001111000000011000000111100000011000110100100;
XPCT = 108'b111000000100000011110000001100110100011001111100001011011111110000101111001111011111110111011111001100111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1000

pattern = 5; // 1000
ALLPIS = 207'b110001011000100011101000001110101110101000011111010111000011100101001101110100111101111001110111001001111001110000110101001011000111000010101110110100000100101100000111100000001100000011110000001100011010010;
XPCT = 108'b111100000110000001111000000100011010110111111111111111111001100000101110010110100110110011000001100010110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1200

pattern = 6; // 1200
ALLPIS = 207'b000010001110101100101000111001010000000101000001000000000000010100010000100001011010001010100100000011011011000110110111111100110111111100000001000000000011101001110101010011000000100110000111101110010001010;
XPCT = 108'b000010010000010011000011110110010001010111111001011010000110100111001111101010001011100110111001110011011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1400

pattern = 7; // 1400
ALLPIS = 207'b000001000111010110010100011100101000000010100000100000000000001010001000010000101101000101010010000001101101100011011011111110011011111110000000100000000001110100111010101001100000010011000011110111001000101;
XPCT = 108'b001101001000001001100001111011001000100101111000101110001111010010001111011111011111110000011001100000001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1600

pattern = 8; // 1600
ALLPIS = 207'b011010000001010110010110110000010011010000011110111011100001100011110010010011010010010100110110100111010001001111000000100110011001100010010110001010000001000101101011110111110110101110011110010011111000001;
XPCT = 108'b001110111011010111001111001011111000011011111011011010011111100110011111101100011000110010111110011001000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1800

pattern = 9; // 1800
ALLPIS = 207'b001101000000101011001011011000001001101000001111011101110000110001111001001001101001001010011011010011101000100111100000010011001100110001001011000101000000100010110101111011111011010111001111001001111100000;
XPCT = 108'b000111011101101011100111100101111100111011111011110100010000010111101110001001000000100101011110111100001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2000

pattern = 10; // 2000
ALLPIS = 207'b100110100000010101100101101100000100110100000111101110111000011000111100100100110100100101001101101001110100010011110000001001100110011000100101100010100000010001011010111101111101101011100111100100111110000;
XPCT = 108'b111111101110110101110011110000111110001101111100000001001111001000011111110100010010111010000001001110011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2200

pattern = 11; // 2200
ALLPIS = 207'b101001110010110111101110001000000101001011001101011100111101101010101000001001011110100100111001010011011101110111010101011101100111010001000100101011010001110111011011111101111000010010001100011010000011011;
XPCT = 108'b111111101100001001000110001110000011111011111100101111010000101011101110111011000110100011111001001011001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2400

pattern = 12; // 2400
ALLPIS = 207'b001110011011100110101011111010000101110100101000000101111111010011100010011111101011100100000011001110001001000101000111110111100111110101110100001111101001000100011011011101111010101110111001100101011101110;
XPCT = 108'b001011101101010111011100110001011101011111111010001010011111110001001111001110100001110010000110110100101110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2600

pattern = 13; // 2600
ALLPIS = 207'b000111001101110011010101111101000010111010010100000010111111101001110001001111110101110010000001100111000100100010100011111011110011111010111010000111110100100010001101101110111101010111011100110010101110111;
XPCT = 108'b000101111110101011101110011010101110011001111000000000001111010001011011001110100010110100000000010000100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2800

pattern = 14; // 2800
ALLPIS = 207'b011001000100000100110110000000100110001100000100101010111110010010001110111100111110001111011111010100000101101111111100100100101101100000001011011001111011101110110000010100011000001100010001110001001011000;
XPCT = 108'b000010100100000110001000111001001011101010111001111110010110101100001111001011011100100111111110111000011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3000

pattern = 15; // 3000
ALLPIS = 207'b001100100010000010011011000000010011000110000010010101011111001001000111011110011111000111101111101010000010110111111110010010010110110000000101101100111101110111011000001010001100000110001000111000100101100;
XPCT = 108'b000001010110000011000100011100100101100011011010101110000000000011010100110011110101100111111110001011110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3200

pattern = 16; // 3200
ALLPIS = 207'b011100110011111100010001011110001110110010001111100001001110000010010101110100001011010101101000010010100110100101010010010000011111000101010100101100011111000100011010100110000000100100111011110100001110101;
XPCT = 108'b001100110000010010011101111000001110100111111011111110011111111100100101010100111100110111011000111111001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3400

pattern = 17; // 3400
ALLPIS = 207'b010100111011000011010100010001000000001000001001011011000110100111111100100001000001011100101011101110110100101100000100010001011011111111111100001100001110011101111011110000000110110101100010010010011011001;
XPCT = 108'b001110000011011010110001001010011011110011111011111110001111110111101011001101111000110100111111001101110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3600

pattern = 18; // 3600
ALLPIS = 207'b001010011101100001101010001000100000000100000100101101100011010011111110010000100000101110010101110111011010010110000010001000101101111111111110000110000111001110111101111000000011011010110001001001001101100;
XPCT = 108'b000111000001101101011000100101001101010011111010000000011111000010011111100100000000111001111111111011001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3800

pattern = 19; // 3800
ALLPIS = 207'b000101001110110000110101000100010000000010000010010110110001101001111111001000010000010111001010111011101101001011000001000100010110111111111111000011000011100111011110111100000001101101011000100100100110110;
XPCT = 108'b001111100000110110101100010000100110100101111000100100000000000110101110101010000010100011011111111010110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4000

pattern = 20; // 4000
ALLPIS = 207'b000010100111011000011010100010001000000001000001001011011000110100111111100100001000001011100101011101110110100101100000100010001011011111111111100001100001110011101111011110000000110110101100010010010011011;
XPCT = 108'b001011110000011011010110001010010011010011111010000000011111111010111111000111110001110100000000000011100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4200

pattern = 21; // 4200
ALLPIS = 207'b000001010011101100001101010001000100000000100000100101101100011010011111110010000100000101110010101110111011010010110000010001000101101111111111110000110000111001110111101111000000011011010110001001001001101;
XPCT = 108'b001101110000001101101011000101001001110010111011111110001111111100011111001101000100110010111111110010110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4400

pattern = 22; // 4400
ALLPIS = 207'b111010001011001011011010010110100101010001011110111001010111101011111001100010000110110100100110110000111010010111110101010001110110101010101001100010011001100011001101010100100110101010010100101100111000101;
XPCT = 108'b110010101011010101001010010100111000010111111111011011001111011111101111100110001001111010011110010000011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4600

pattern = 23; // 4600
ALLPIS = 207'b100111100111011000110001110101010101111001100001110111001010010011001010101010000111101100001100111111111010110101010111110001101111001000000010101011001101001110010000001001010101110010110101111110000000001;
XPCT = 108'b110001000010111001011010111110000000001101111111011011111111001001101111001111010110110100011001001101010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4800

pattern = 24; // 4800
ALLPIS = 207'b001001010001010001000100000100101101101101111110010000000100101111010011001110000111000000011001111000011010100100000110100001100011111001010111001111100111011000111110100111101100011110100101010111011100011;
XPCT = 108'b001100111110001111010010101011011100100101011000101110011111111000101111100101000100111010100000011100110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5000

pattern = 25; // 5000
ALLPIS = 207'b100100101000101000100010000010010110110110111111001000000010010111101001100111000011100000001100111100001101010010000011010000110001111100101011100111110011101100011111010011110110001111010010101011101110001;
XPCT = 108'b111010011011000111101001010111101110111001111100101111011111001000101111100101111011110011100000010100110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5200

pattern = 26; // 5200
ALLPIS = 207'b001000110110101001001101111111001100001010010001001111100000101101000010101000100101000110011001111001100001010111101100110001001100100011000011101001111000001001111001001010111101100000010110111101101011011;
XPCT = 108'b000001011110110000001011011101101011111111111010101110000000010000000100101011000101101101111000110111010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5400

pattern = 27; // 5400
ALLPIS = 207'b100100011011010100100110111111100110000101001000100111110000010110100001010100010010100011001100111100110000101011110110011000100110010001100001110100111100000100111100100101011110110000001011011110110101101;
XPCT = 108'b110100100111011000000101101110110101101101111110101111001111011100111111111100101100111100011110011001010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5600

pattern = 28; // 5600
ALLPIS = 207'b101000101111010111001111100001110100010011101010111000011001101101100110110001001101100111111001111001111111101011010110010101000111010101100110100000011111111101101000110001101001111111111010000111000110101;
XPCT = 108'b110110001100111111111101000011000110100111111100101111011111110100111111111100001010110000111110011100100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5800

pattern = 29; // 5800
ALLPIS = 207'b010100010111101011100111110000111010001001110101011100001100110110110011011000100110110011111100111100111111110101101011001010100011101010110011010000001111111110110100011000110100111111111101000011100011010;
XPCT = 108'b000011001010011111111110100011100011101011101001111110011111001010110101011101110011110000111110100011100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6000

pattern = 30; // 6000
ALLPIS = 207'b101010001011110101110011111000011101000100111010101110000110011011011001101100010011011001111110011110011111111010110101100101010001110101011001101000000111111111011010001100011010011111111110100001110001101;
XPCT = 108'b111001100101001111111111010001110001001001101100001011101111101001011111111110000111110001111110111110001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6200

pattern = 31; // 6200
ALLPIS = 207'b110101000101111010111001111100001110100010011101010111000011001101101100110110001001101100111111001111001111111101011010110010101000111010101100110100000011111111101101000110001101001111111111010000111000110;
XPCT = 108'b110000110110100111111111101000111000110011101111111111101111000001001111011111100111111011100001000000111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6400

pattern = 32; // 6400
ALLPIS = 207'b101011011010010100110011110000101111010110011100011101000100100101000110010001101101111100100000101000111010001010111001001100100001010111010001011011011100010001100100001011010101110111011100010011111011001;
XPCT = 108'b110001010010111011101110001011111011001001111111011011111001001010001110010100100010111011100001011011111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6600

pattern = 33; // 6600
ALLPIS = 207'b100011011001100011111110011001001001000111110110110100101011011000101111101011101101000111010001000101101001010000101110111111010010000101001010011011010110101011111010010011000001010101010110101110001011111;
XPCT = 108'b111010010000101010101011010110001011000111111100001011001111000101011111000101010000110100000111010110000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6800

pattern = 34; // 6800
ALLPIS = 207'b100111011000011000011000101101111010001111000011100000011100100110011011010110101101011010101001110011000000111101100101000110101011101100000111111011010011110110110101011111001011000100010011110000110011100;
XPCT = 108'b110011110101100010001001111000110011010011111101011011100000010000000110000000000100100010011111111001000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7000

pattern = 35; // 7000
ALLPIS = 207'b000101011000100101101011110111100011101011011001001010000111011001000001001000001101010100010101101000010100001011000000111010010111011000100001001011010001011000010010111001001110001100110001011111101111101;
XPCT = 108'b001111000111000110011000101111101111100111111001111110000000010110111110010001100100100100011110011010101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7200

pattern = 36; // 7200
ALLPIS = 207'b010111100010100000111101011100100110010110001110101000101000111100011100110001011000101100000100001011110001010111000010010111100111011000101010100100001100110101001100111000111000001101110100110000001101100;
XPCT = 108'b000111001100000110111010011000001101001011111001011010000000101001101110011001100100101001011110100111111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7400

pattern = 37; // 7400
ALLPIS = 207'b001011110001010000011110101110010011001011000111010100010100011110001110011000101100010110000010000101111000101011100001001011110011101100010101010010000110011010100110011100011100000110111010011000000110110;
XPCT = 108'b001011100110000011011101001100000110001011111001011010001111001100001111101110000101111010000110010111110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7600

pattern = 38; // 7600
ALLPIS = 207'b110011001100000001101000110110010111001001011011010000000011000101001011101111001101110010000000010011001000000000000010111100111011011000101000011111111011101110011011011000100101101101100101101011110101000;
XPCT = 108'b111011001010110110110010110111110101010011111101011011010000010010001110000000110101101111111110000011111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7800

pattern = 39; // 7800
ALLPIS = 207'b111001100110000000110100011011001011100100101101101000000001100010100101110111100110111001000000001001100100000000000001011110011101101100010100001111111101110111001101101100010010110110110010110101111010100;
XPCT = 108'b110101100001011011011001011001111010111111111101111111100000010010101100000000011000100011011110000101100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8000

pattern = 40; // 8000
ALLPIS = 207'b011100110011000000011010001101100101110010010110110100000000110001010010111011110011011100100000000100110010000000000000101111001110110110001010000111111110111011100110110110001001011011011001011010111101010;
XPCT = 108'b001110110100101101101100101110111101100011111001111110000110111111101111010001111010101001011110101110100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8200

pattern = 41; // 8200
ALLPIS = 207'b011000101101001001101010100111101100010101110011100000001001010010100101111110100010010111010001010011101101010101110010001110100101110101100111110101000111111110111011001101101111000011010100001010101000110;
XPCT = 108'b001001101111100001101010000110101000110011010001111110011111101000011111100111000111111110111000011100111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8400

pattern = 42; // 8400
ALLPIS = 207'b111010100010001101010010110010101000100110000001001010001101100011011110011100001010110010101001111000000010111111001011011110010000010100010001001100011011011100010101110000011100001111010010100010100010000;
XPCT = 108'b110110000110000111101001010010100010011011110101011011001111100111101111101110011010110011100000011000101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8600

pattern = 43; // 8600
ALLPIS = 207'b111000011100001010110011001101110100100101011000101000101010010010111011000100011001010101101011001111110100111010000000101110100110101011100110100101111110010100001101001010101100101101001100001111011110111;
XPCT = 108'b110001011110010110100110000111011110110111111101111111010000011000011110000010110111100010011001110001011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8800

pattern = 44; // 8800
ALLPIS = 207'b011100001110000101011001100110111010010010101100010100010101001001011101100010001100101010110101100111111010011101000000010111010011010101110011010010111111001010000110100101010110010110100110000111101111011;
XPCT = 108'b001100100011001011010011000011101111101111111001111110010000011101111110110000001110100110111001110011100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9000

pattern = 45; // 9000
ALLPIS = 207'b011000110011101011001011010010000011100101101110110000000011101110100010010010011101101100011011100010001001011011010010010010101011000100011011011111100111000110001011000100000000100101101011100100000001110;
XPCT = 108'b001000100000010010110101110000000001110111111001111110001111000111111111100101111111110110011001101100110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9200

pattern = 46; // 9200
ALLPIS = 207'b111010101101011100000010001000011111011110001111100010001000111101011101101010010101001111001100100000110000111000011011010000010111001100101111011001001011000000001101110100101011111100001101010101110110100;
XPCT = 108'b110110101101111110000110101001110110010111111101011011101111000110111111000100101010110000111111101111101110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9400

pattern = 47; // 9400
ALLPIS = 207'b111101010110101110000001000100001111101111000111110001000100011110101110110101001010100111100110010000011000011100001101101000001011100110010111101100100101100000000110111010010101111110000110101010111011010;
XPCT = 108'b111111010010111111000011010110111011101011111111111111010000011100001100110001110000100000000111111000011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9600

pattern = 48; // 9600
ALLPIS = 207'b011110101011010111000000100010000111110111100011111000100010001111010111011010100101010011110011001000001100001110000110110100000101110011001011110110010010110000000011011101001010111111000011010101011101101;
XPCT = 108'b001011100101011111100001101001011101010111111001011010011111010011001111100111010011110000011001100100110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9800

pattern = 49; // 9800
ALLPIS = 207'b100111101010110101110000001000100001111101111000111110001000100011110101110110101001010100111100110010000011000011100001101101000001011100110010111101100100101100000000110111010010101111110000110101010111011;
XPCT = 108'b110110110001010111111000011001010111001101111101010001010000100001101100010001001101101101000000010110111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10000

pattern = 50; // 10000
ALLPIS = 207'b100101000001110011011111100101001110010010000100100101001101011011110110011000001111010011011111001000110101110100000010101111100010000000111011101000001010110101001000001101000010111001000000111101011101110;
XPCT = 108'b110001100001011100100000011101011101100111110110100101001111010111111111110110111000111001100111101001010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10200

pattern = 51; // 10200
ALLPIS = 207'b100100010100010000001000010011111001100101111010101000101111100111110111101111011100010000101110110101101110101111110011001110110011101110111111000010111101111001101100010000001010110010011000111001011000100;
XPCT = 108'b110010000101011001001100011101011000100011111100100101001111110010101111111101101011111100100000110100001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10400

pattern = 52; // 10400
ALLPIS = 207'b100100111110100001100011101000100010011110000101101110011110111001110111010100110101110001010110001011000011000010001011111110011011011001111101010111100110011111111110011110101110110111110100111011011010001;
XPCT = 108'b111011111111011011111010011111011010100001011100100101011111001111011111110100110011110100000001010110110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10600

pattern = 53; // 10600
ALLPIS = 207'b110010011111010000110001110100010001001111000010110111001111011100111011101010011010111000101011000101100001100001000101111111001101101100111110101011110011001111111111001111010111011011111010011101101101000;
XPCT = 108'b111001110011101101111101001101101101011111111111011011101111001100111111101111110101111000011110000100011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10800

pattern = 54; // 10800
ALLPIS = 207'b101111111011000001111111011011010110001011011001100001101110100100010001010110010110100101010100110011000100100101010000100110100100011000111101100011000001000100110111110001000000000011000101101001000000111;
XPCT = 108'b111110000000000001100010110101000000010011111111011011001111110011010111011101101000110000011000001011010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11000

pattern = 55; // 11000
ALLPIS = 207'b110111111101100000111111101101101011000101101100110000110111010010001000101011001011010010101010011001100010010010101000010011010010001100011110110001100000100010011011111000100000000001100010110100100000011;
XPCT = 108'b111111001000000000110001011000100000010111111101011011011001000001011100111110110011111100111001100101011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11200

pattern = 56; // 11200
ALLPIS = 207'b110110100101001100111100001011110101100111000111010001001001010001100100011011011111001000001010001110100010101110010011001000010101110100010110110111000100011001000010110101011101110111000100111110110011001;
XPCT = 108'b111110100110111011100010011110110011001111111111011011101111101101001111110111011000110011111111100000111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11400

pattern = 57; // 11400
ALLPIS = 207'b011011010010100110011110000101111010110011100011101000100100101000110010001101101111100100000101000111010001010111001001100100001010111010001011011011100010001100100001011010101110111011100010011111011001100;
XPCT = 108'b000011011111011101110001001111011001010111111001011010000000101111111110111010001011101111111111111001111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11600

pattern = 58; // 11600
ALLPIS = 207'b101101101001010011001111000010111101011001110001110100010010010100011001000110110111110010000010100011101000101011100100110010000101011101000101101101110001000110010000101101010111011101110001001111101100110;
XPCT = 108'b110101100011101110111000100111101100101111111101111111001111001100101111111110000110110001100110101001101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11800

pattern = 59; // 11800
ALLPIS = 207'b100101111010100111110011010000001100101111100011001100010011111001011001001110111100111101010100111001000101011001010100010001011101001100010011111010100011000111111001110000011010010001001011100001010101001;
XPCT = 108'b110110000101001000100101110001010101111001111100101111110110001001011111010001111011101001011110000010101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12000

pattern = 60; // 12000
ALLPIS = 207'b111001001000011100011111001000011111001000110111111110101110001110011110111010100111100100000011101110101000011110000010101010010100111110101110001000010111101100001111011000111001101010110010110010000000111;
XPCT = 108'b111011001100110101011001011010000000111011111101111111000000100100010110001011101110100100111110111100010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12200

pattern = 61; // 12200
ALLPIS = 207'b110111010001000001101001000100010110111011011101100111110000110101111101000000101010001000101000000101011110111101101001110111110000000111110000110001001101111001110100001100101000010111001110011011101010000;
XPCT = 108'b110001101100001011100111001111101010000011101111011011111111110011010111111110000100111000111111001110101110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12400

pattern = 62; // 12400
ALLPIS = 207'b101000001110110111101001000001001001000001010100010101101111110100000110011110110110011111011110111000010010110110001110001100100001001101101111110110110000011001100100110011010000010100111000000111101111101;
XPCT = 108'b110110010000001010011100000011101111101111111111111111111111101010110101011110001000110101000001011111101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12600

pattern = 63; // 12600
ALLPIS = 207'b001100001001101010100010000000010110000000111101011100000011110000111110001001010001010111111000011001101010001000110011011011110000110111000011110110100001101111000011111110100011101000010101110010111101000;
XPCT = 108'b001111111001110100001010111010111101110001111001110100001111011110010101100110000010111010011001110010011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12800

pattern = 64; // 12800
ALLPIS = 207'b000110000100110101010001000000001011000000011110101110000001111000011111000100101000101011111100001100110101000100011001101101111000011011100001111011010000110111100001111111010001110100001010111001011110100;
XPCT = 108'b000111110000111010000101011101011110011001111001011010011111010010111011000101100010110100000001011111000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13000

pattern = 65; // 13000
ALLPIS = 207'b001010010100000010110010110000011011101111000001110011000111101100110101101100110011110000010110110001000111100011101110111001100100011110011111101011110010000010001011111111000000111111010101101100111101110;
XPCT = 108'b001111110000011111101010110100111101010101111010000000010000111111011010001010110000100000000111001011000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13200

pattern = 66; // 13200
ALLPIS = 207'b001110111111001110111111111000010100101000100110100001000100000100101000101011100000000010100010101010101001000011011111111110001000010111101000000000111111001110110110011111010100111101111101110100110100100;
XPCT = 108'b001011110010011110111110111000110100001111111011011010011111011101011111011100100001110001011001011010010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13400

pattern = 67; // 13400
ALLPIS = 207'b000111011111100111011111111100001010010100010011010000100010000010010100010101110000000001010001010101010100100001101111111111000100001011110100000000011111100111011011001111101010011110111110111010011010010;
XPCT = 108'b001001111101001111011111011110011010010011111000001010011111011100001111101110100110111000000000111101011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13600

pattern = 68; // 13600
ALLPIS = 207'b001000011010111100001001011110011100010101001111110000110110110011111000010111000001111010000001011000100000100010011111011101011000011101011101110101001001111100011110000111000001101101001000011111100111010;
XPCT = 108'b001000110000110110100100001111100111100111111000100100010110111010101111111000111111100010100110010011111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13800

pattern = 69; // 13800
ALLPIS = 207'b100100001101011110000100101111001110001010100111111000011011011001111100001011100000111101000000101100010000010001001111101110101100001110101110111010100100111110001111000011100000110110100100001111110011101;
XPCT = 108'b111000011000011011010010000111110011110101111100100101101111100000001111001111011111110100011110000001011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14000

pattern = 70; // 14000
ALLPIS = 207'b010111001100111111110100111011100110010010001100101010110010111101110100010001111101001000101101000000001011101111101111001000001100010111011111100001001100000111101001100000010110111110110101100000000011101;
XPCT = 108'b000100000011011111011010110000000011011011111001011010001111110010011111101101101011111000000000001001010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14200

pattern = 71; // 14200
ALLPIS = 207'b000101110011001111111101001110111001100100100011001010101100101111011101000100011111010010001011010000000010111011111011110010000011000101110111111000010011000001111010011000000101101111101101011000000000111;
XPCT = 108'b001011000010110111110110101100000000100011111000101110001001010000011010011101011010110100011001000111101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14400

pattern = 72; // 14400
ALLPIS = 207'b100011011011010110011001001001101110010011100010000001110010010111001001110101011010000000111000101000001010100101110111111100101010000000001001001010000100010111111100110011110100001111101010101001101010011;
XPCT = 108'b110110011010000111110101010101101010001011111110001011011111000111001101011101111000111001000000100111101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14600

pattern = 73; // 14600
ALLPIS = 207'b000110111001011101110011100010001110010100011101110100101000101110011001001110010011100111110011000001001101000010100001001100101101110100110110011101000100001101110101011100010011110000100110001001100101110;
XPCT = 108'b000011100001111000010011000101100101011001011001011010001111111011000101000100010011111100011001000101000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14800

pattern = 74; // 14800
ALLPIS = 207'b100011011100101110111001110001000111001010001110111010010100010111001100100111001001110011111001100000100110100001010000100110010110111010011011001110100010000110111010101110001001111000010011000100110010111;
XPCT = 108'b111101110100111100001001100000110010000111111100001011000000010001011110011000000000100101000110010100011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15000

pattern = 75; // 15000
ALLPIS = 207'b101101001101101100011101001100011101011101000000100010110110111100101010000111001110100001101010100001001100110001000000011000111000100010110101001001001011100110010111011011111000001111001111010000011001100;
XPCT = 108'b111011011100000111100111101000011001111011111101111111001111101000101011000101000011110100011000001101110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15200

pattern = 76; // 15200
ALLPIS = 207'b111101010011111001101000000110010111110001100110001001111100101100100111011110011110101010011100100010101100101010001000101110100110001001111101010001100011111100111000001101001000100101110000101010100110101;
XPCT = 108'b110001100100010010111000010110100110100011111111111111101111100110111111011101010101110111111001100111001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15400

pattern = 77; // 15400
ALLPIS = 207'b011110101001111100110100000011001011111000110011000100111110010110010011101111001111010101001110010001010110010101000100010111010011000100111110101000110001111110011100000110100100010010111000010101010011010;
XPCT = 108'b000000111010001001011100001001010011000111111001011010000110111001011111010000001111101110011111110111100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15600

pattern = 78; // 15600
ALLPIS = 207'b101111010100111110011010000001100101111100011001100010011111001011001001110111100111101010100111001000101011001010100010001011101001100010011111010100011000111111001110000011010010001001011100001010101001101;
XPCT = 108'b111000010001000100101110000110101001001011111100001011100000000100111110111000101111101100111111111001110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15800

pattern = 79; // 15800
ALLPIS = 207'b010111101010011111001101000000110010111110001100110001001111100101100100111011110011110101010011100100010101100101010001000101110100110001001111101010001100011111100111000001101001000100101110000101010100110;
XPCT = 108'b001000001100100010010111000001010100010111111011011010001111001000001111101110100010110110000000000110000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16000

pattern = 80; // 16000
ALLPIS = 207'b010101100010100111100110100011110101111000010001011110011111000101001110101110110100110010001001110000111101001100101111010101101100011000011100100100011111011001100000010011001010000110000101101101100001101;
XPCT = 108'b000010010101000011000010110101100001100111011001111110000000000101111110000011111101100010011111110100100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16200

pattern = 81; // 16200
ALLPIS = 207'b100101111111100000101001000110010001101011011011111010100011011111000000001100011000001101011100000110100100000011011101000101110111110111010001010010110011001110011100011000110110010101110111110110111101010;
XPCT = 108'b110011001011001010111011111010111101101111111100101111111111001011011111101100010001110111011110100100100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16400

pattern = 82; // 16400
ALLPIS = 207'b100011101110101011111001000000011110100110111110010001100111010101010111010100011100011010010011111001110111100110100000111011101011110001111010000110100011011111010111001111101000100110011111001011011111100;
XPCT = 108'b111001111100010011001111100111011111010011110111011011100000000110101110110010101100101000111111011100010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16600

pattern = 83; // 16600
ALLPIS = 207'b110010001010111001001101000001111101010101100111001011010110010111110010100010011101011111100000000110000011011111111111100100001100110000010000110011100111011011000101111010011111001010100101000100000111001;
XPCT = 108'b110111010111100101010010100000000111011111111111011011101111000001010101100110000000111010000001001101111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16800

pattern = 84; // 16800
ALLPIS = 207'b000110010011111101100000000001100101101001010001011101111010000111011011111111111101001110111100111001111110010001101000010011110101000000001010011110110110011010000001010111000010110001101011100111110001000;
XPCT = 108'b000010110001011000110101110011110001010101111011011010011111110001111111100110101001111100111111011010001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17000

pattern = 85; // 17000
ALLPIS = 207'b000011001001111110110000000000110010110100101000101110111101000011101101111111111110100111011110011100111111001000110100001001111010100000000101001111011011001101000000101011100001011000110101110011111000100;
XPCT = 108'b000101011000101100011010111011111000000001111001011010001111001011101111111101100111111001111001111001000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17200

pattern = 86; // 17200
ALLPIS = 207'b010100000110011000111110100011101100100010000101001001000001100100111000010001001011100001100110111110100010101000110101010001010001001000011110000011110010111111000000000110111010101010011111010100011101111;
XPCT = 108'b000000111101010101001111101000011101101111111011111110000000001010001110111001101101101010000110000000000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17400

pattern = 87; // 17400
ALLPIS = 207'b110001000100001000110000101100000000101000110000000110010011001011000000001111000000111010100000000110001100101110000111110111000011001101101010100011001110110111100000010110111001111010101000011110100111001;
XPCT = 108'b110010111100111101010100001110100111101111111101111111111111000100111111100101100010110100000001110101110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17600

pattern = 88; // 17600
ALLPIS = 207'b110110100000010001111111011010111010110110000100101110101011010000010111010100101010010111101100111001111101101101110110010111000110111111010100111010111100000001001000001100001011011101101000110001011001000;
XPCT = 108'b110001100101101110110100011001011001000011011101011011001111011011001111110111010111110000000000111011011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17800

pattern = 89; // 17800
ALLPIS = 207'b011011010000001000111111101101011101011011000010010111010101101000001011101010010101001011110110011100111110110110111011001011100011011111101010011101011110000000100100000110000101101110110100011000101100100;
XPCT = 108'b000000110010110111011010001100101100000011101011011010001111010111111111111110111011111011000001001011001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18000

pattern = 90; // 18000
ALLPIS = 207'b010110001010011110011010001111010111100001000101111001111100010100111010111011010011001000100111000011110100110010111101010110110001100001110010010001111101100110000001001100101000011000010110110110000110100;
XPCT = 108'b000001101100001100001011011010000110010111111011011010001111011101101111100110110101111001100001001011111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18200

pattern = 91; // 18200
ALLPIS = 207'b101011000101001111001101000111101011110000100010111100111110001010011101011101101001100100010011100001111010011001011110101011011000110000111001001000111110110011000000100110010100001100001011011011000011010;
XPCT = 108'b110100110010000110000101101111000011001011111101011011011111111011111111100101100010111010000000101100000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18400

pattern = 92; // 18400
ALLPIS = 207'b001001010001100010110111100111100000001110011011001011110010011000000000110111100011101111001011011101110111011110010001110011111100011100010000110100000011011100000100111100010100100010110110110100011101111;
XPCT = 108'b000111100010010001011011011000011101101101111011111110001111000100001011000100000010111101100111011011101001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18600

pattern = 93; // 18600
ALLPIS = 207'b011011000101111010011010011110011000001101111101111001001110111110000000111010011011010100111001101010101010101001110101101111000011011011010100111001000011101011000101110011010001101010011011011001011010100;
XPCT = 108'b000110010000110101001101101101011010011011111011011010001111010100111111111100100101110100011111111110100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18800

pattern = 94; // 18800
ALLPIS = 207'b001011001000001101001010110011110110001010001001110000011000111011100000100010110100101101100000101001100110011011000100010001110010100100101101100000010010001000110111111110101010101001001011011000000101101;
XPCT = 108'b001111111101010100100101101100000101010011111001011010000000010011010010101011100101100101011110000110011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19000

pattern = 95; // 19000
ALLPIS = 207'b001011100011100001100101001011011101101100111001010111110100010110111000111111001110100100010011010111101110111000100000110111100000110101011011101100000111111110001001000011111110001000100100000010011100100;
XPCT = 108'b000000011111000100010010000010011100011001101010000000001111010111111111000101110011111000111110011101111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19200

pattern = 96; // 19200
ALLPIS = 207'b100101110001110000110010100101101110110110011100101011111010001011011100011111100111010010001001101011110111011100010000011011110000011010101101110110000011111111000100100001111111000100010010000001001110010;
XPCT = 108'b110100001111100010001001000001001110101001110111111111011111110011101111000110000111110101111110100000000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19400

pattern = 97; // 19400
ALLPIS = 207'b111101110100101101010111011010101011101010101010101111000111101110110111011100001000000011000111110100000110011000001100111111000010001000100011000111100001010001110011010110010101100000011111111010011101011;
XPCT = 108'b111010110010110000001111111110011101111011111111111111010000001001011110000001101001101110100001101000001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19600

pattern = 98; // 19600
ALLPIS = 207'b100011110100011111010110001100010001011011011011110101001110100010011101010010011111011001000110111110101100011110110111111000100010111100100111111001101100110010000110110010011111100101001101010000001101110;
XPCT = 108'b111110010111110010100110101000001101001001111111011011100000011010001010101011111011101111100111000010001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19800

pattern = 99; // 19800
ALLPIS = 207'b110001100111110000010110100101110010000010001101110000100010100000010011000110000001100011100110000100111001010010101111110101000110000101111100010001001111010100010110010100001101001111000100000100010010101;
XPCT = 108'b111010100110100111100010000000010010100111111101111111001111110011001011111101010010111011011111001110011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20000

pattern = 100; // 20000
ALLPIS = 207'b110100100100111100111001111110001110100010100111011101010001100000110100111101100001110111110000000000000011101000110100110011101101100001110111010011010001110100101111100101110000111101101111001100001000011;
XPCT = 108'b111100101000011110110111100100001000111111111111111111010110011001001111001010011100100000111111010010111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20200

pattern = 101; // 20200
ALLPIS = 207'b111010010010011110011100111111000111010001010011101110101000110000011010011110110000111011111000000000000001110100011010011001110110110000111011101001101000111010010111110010111000011110110111100110000100001;
XPCT = 108'b111110011100001111011011110010000100011111111101011011111111111000001111101110101010110001000001000101111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20400

pattern = 102; // 20400
ALLPIS = 207'b100101000110001011011110011110000000111001101100101111001001100000000011011110001110111100101101110111011101111001000111001111110001110001000011010000001101110000010011110001010010001011011011010001110111111;
XPCT = 108'b111110000001000101101101101001110111111011111111111111100000101010111110100010011101100100111110001111010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20600

pattern = 103; // 20600
ALLPIS = 207'b101100000001011100000100001011001010111111001011011000110010110000111001011111010111101001011000010010010101011000110110010010011111001001100001000001010011111111001101111111001111110110100110001111111111111;
XPCT = 108'b110111110111111011010011000111111111110101111100100101100110011111101111100001100010100100111111011110010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20800

pattern = 104; // 20800
ALLPIS = 207'b101100110110011110100001111101001100110011100011001001110001011001100001010001000010101011010011100000011001001010000110100010000011111100000110010111101110101000000010101111100100100000111110010010000101111;
XPCT = 108'b111101111010010000011111001010000101100001111111111111100000011101111110011000000100101111000001100010111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21000

pattern = 105; // 21000
ALLPIS = 207'b010101011100001000110100010101101111110101010100100100011010000111001111110110101011100010110001010100111011001011010111010100001111001000010100111001010011010110001001100010101101010011000001001001111011101;
XPCT = 108'b000100011110101001100000100101111011110011111001111110000110011010111011110011111111100111011111011010110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21200

pattern = 106; // 21200
ALLPIS = 207'b110111100101110011101001011010011110110111100001110011001100010010001011011010100111100000100010100000001001011000101110110000110011101011111010101011101101110001111001000011010111111001100011100101110001100;
XPCT = 108'b110000010011111100110001110001110001011111111111011011001111000000001011000110011101110010011111101000100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21400

pattern = 107; // 21400
ALLPIS = 207'b111011110010111001110100101101001111011011110000111001100110001001000101101101010011110000010001010000000100101100010111011000011001110101111101010101110110111000111100100001101011111100110001110010111000110;
XPCT = 108'b110100001101111110011000111010111000000011010111011011001001010111011110100101100100110101000001000001100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21600

pattern = 108; // 21600
ALLPIS = 207'b010111011110010111001110100101101001111011011110000111001100110001001000101101101010011110000010001010000000100101100010111011000011001110101111101010101110110111000111100100001101011111100110001110010111000;
XPCT = 108'b001100100110101111110011000110010111010111111011011010011001110110011110100111110110110111000000001000011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21800

pattern = 109; // 21800
ALLPIS = 207'b010111000101010100010111110110011111010100000011011011111001111111101010101100010111111111101110010111100111100011000011101011000000101010010100011111010010101001101010100010111111111010101010010100001010101;
XPCT = 108'b001100011111111101010101001000001010001111111011011010001111010000011111101101110110111001111111110110011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22000

pattern = 110; // 22000
ALLPIS = 207'b011011100000111010011001110111011011001100101100100000111000001110101101001001111110110111111110001001000100100001000110000110011111111101110000011011011100010110010011100001111011100101100100001000011000011;
XPCT = 108'b001100001101110010110010000100011000011011111001011010011001110000001000011100010101111110000000011000010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22200

pattern = 111; // 22200
ALLPIS = 207'b101000101001100001111010010111001010001010100111011110001000010010111100110000100100100101111010001110101100010001100111011101001000001000001001011010011111111001101101110001001010100010010111101111011100110;
XPCT = 108'b110110000101010001001011110111011100110111111100100101011111001100111111101110001010111110011111000010001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22400

pattern = 112; // 22400
ALLPIS = 207'b100101011010100010111111000101111010101100101010001101101000001001100100001011000101011100011011011100011001000001000100110111111000110101110100101011110010101001100010100110100000101110100001000010101010101;
XPCT = 108'b111100111000010111010000100010101010100011111111111111101111100010000111000101010100111111000000110110110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22600

pattern = 113; // 22600
ALLPIS = 207'b000111110011011010001000010110101101001101010010110100011111010000101011000111111100111111110011000111001101110000000001001000101101000111101101100001110110010100000111100100001010111001010001110010001101100;
XPCT = 108'b001100100101011100101000111010001101010011111001011010001111001010111111110101101100111000011110000101110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22800

pattern = 114; // 22800
ALLPIS = 207'b000101010100100010011101101110101010000101000010101011101010110101111101000010011001100100100011101011001001100011101011010100110001000010111000110101101011001011101101000100111101010110011010011000011011011;
XPCT = 108'b000000101110101011001101001100011011111011111010100100010000010000111010001011011000101110111111101010110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23000

pattern = 115; // 23000
ALLPIS = 207'b101111010000100101011011101011001011011111100111010010101000010011001100000101001011011011101110001011001010101001010101111110110000100101001001110000101001001000011010011111100001110110100110101110111010010;
XPCT = 108'b111011111000111011010011010110111010000111111100001011110000111011101010010010110011100100100000010000110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23200

pattern = 116; // 23200
ALLPIS = 207'b001100001010010000110100100100000111100000101110110010001011111101001001110100001011011101101011011111010001010101111010000110111000101001100001001110000011111010001111001000100101001001010010000000000000111;
XPCT = 108'b001001001010100100101001000000000000110001111000101110010000011001000100100011000111101011111110110000110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23400

pattern = 117; // 23400
ALLPIS = 207'b110111000100000100110010100011000100011110111010110110111111101001011111101101011101100000111000110101101000000010100001110011000001110110001011101100101110111100000100001110101011100100000010101110111011101;
XPCT = 108'b110001111101110010000001010110111011000111111101011011001001110001101110100100000000111100000001111000001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23600

pattern = 118; // 23600
ALLPIS = 207'b111100000010111110011001001111011001110010110100011101110010010110001001000111010111011110100000110000000010001011000000101011011001110110101001000111011000100000101011011011110100101101101010010101111000001;
XPCT = 108'b111011011010010110110101001001111000111111111111111111110000101001001110101000110001100011011111101101100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23800

pattern = 119; // 23800
ALLPIS = 207'b011110000001011111001100100111101100111001011010001110111001001011000100100011101011101111010000011000000001000101100000010101101100111011010100100011101100010000010101101101111010010110110101001010111100000;
XPCT = 108'b000101101101001011011010100110111100011011111001011010011111110010001011001111000110110101011000000100110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24000

pattern = 120; // 24000
ALLPIS = 207'b010011000010010001111111011100101111101110011001011010101110110011101011010110100010101001001000111100000010101001110000100001101111101011000011010110101110101000100001101101001001100110110000110000100110001;
XPCT = 108'b000101100100110011011000011000100110010011111001011010011111010011101111001110010011110000100000001011111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24200

pattern = 121; // 24200
ALLPIS = 207'b011011011001100010100101001111111111011000000100000010110000011000111011101000101010001101110001010011100001110010011110011011010111011011100110101000101111101101011011010110101110010001011001101001100110110;
XPCT = 108'b001010111111001000101100110101100110010011111001011010001111011110001011111100111001110000000000010010000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24400

pattern = 122; // 24400
ALLPIS = 207'b110000001100101110110101111010101000001010101100111101011100011000010110000101110011111100010011011011001111010011110001101001011010101000001111110001110101101010100101011011111110001010011101111110110101011;
XPCT = 108'b110011011111000101001110111110110101111111111111111111100110001110010101001000010001101011111000001110011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24600

pattern = 123; // 24600
ALLPIS = 207'b000011010010011001101101010000110001101110110010110101111100110000010011101011110011100011110001110111001111000010100011011010100000010010100000100111000101000001010111000100111100100010011000000011100101000;
XPCT = 108'b001000101110010001001100000011100101011011111011011010011111101000111111110111110111111101000000000100011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24800

pattern = 124; // 24800
ALLPIS = 207'b100101111001101001111100010000010111110000111111000111111100001110010101000110110010000011111110000000010101000000010100001001010101100101010110110101110001010100101011011010000111111000010011011001010000011;
XPCT = 108'b111011010011111100001001101101010000110011111110101111011111000110101111001101000111110011100001010101000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25000

pattern = 125; // 25000
ALLPIS = 207'b011000101100011101001000000001111000001001001001110010001011011011101010000100100001010000101110010000100011100010000010111000001000011100011100101000010010110001101011101111011111111011101101011111111111000;
XPCT = 108'b001101110111111101110110101111111111111111111001111110001111111110001111000111000110110111100001110111001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25200

pattern = 126; // 25200
ALLPIS = 207'b001010110111001001111110010001001100010101110000000001000010110001001001111011110001000011101010111101100000101001010100010000001001001110101000100100111100000110101000010100101100001000001101101000001110000;
XPCT = 108'b000010101110000100000110110100001110000011111010001010011111100110101011111110111001111011011111000010000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25400

pattern = 127; // 25400
ALLPIS = 207'b100101101100001110111111011010110111001000101100100100100101101010110001110101001111011111011011100111101101110001010110001100100001001100100001100001011011011001011010101101100110111111111110010010000110101;
XPCT = 108'b111101101011011111111111001010000110100010111100100101100110101000111111010010011000100101011110000000011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25600

pattern = 128; // 25600
ALLPIS = 207'b010111000100010110110011110110001011101001000010100011101111111111000111110010001010000010001111100010110010000010001011011010010010011010000101001000010110000110000011011111000101100011101000010110110001001;
XPCT = 108'b001011110010110001110100001010110001010111111011011010010000000000001010110011111001100110111111010101100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25800

pattern = 129; // 25800
ALLPIS = 207'b000100000010010000110101111100010110100111001101010110100000010101100000101101000001000011111010010101001101110000110110100011111101101001010111110011010011101011001110100001111010110010001000010111010100101;
XPCT = 108'b001100001101011001000100001011010100101101111000101110001111010001011111110100101110111100000000111111011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26000

pattern = 130; // 26000
ALLPIS = 207'b101011010011011111000011110000000111100110101100001011010011110100011001000011000011111110001001100101111100100011010110010101010101111001000101011001111101000111111100100100001100011111001011001001101100100;
XPCT = 108'b110100100110001111100101100101101100000001111110001011101111001100011011001100000001111110011110011001000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26200

pattern = 131; // 26200
ALLPIS = 207'b010001001011111000001000100000001100110111000010010101100010000110000101011000111011000110001101000000100001110011011000101110110100010101110011011111010010001110111000010010000000011100111011101100000010000;
XPCT = 108'b000010010000001110011101110100000010100110111011111110011111011000011111111110110000110101111111110100110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26400

pattern = 132; // 26400
ALLPIS = 207'b101000100101111100000100010000000110011011100001001010110001000011000010101100011101100011000110100000010000111001101100010111011010001010111001101111101001000111011100001001000000001110011101110110000001000;
XPCT = 108'b110001000000000111001110111010000001100101111100101111001111111001001111010110000111110011011110111111001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26600

pattern = 133; // 26600
ALLPIS = 207'b010101110100001000010111110100010100011001100110100101000001000011100000011010111111010011001101011011100111111110111101010101110000100010100000001111010000011010010000010110100101001010000111000001110011110;
XPCT = 108'b000010111010100101000011100001110011100010101011111110000000001011101110010001010100100111100110000010000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26800

pattern = 134; // 26800
ALLPIS = 207'b010001111110101000001111111111101000011001011010101001111010100010000110100000110000010000001111110011100001001010100100001000001011101001100110101011010100111010110001000010100001111000111110010000100100101;
XPCT = 108'b000000011000111100011111001000100100110011111011111110001001101110011110011110000011111011100000110100010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27000

pattern = 135; // 27000
ALLPIS = 207'b001000110101011000001111100010110111011100010101001010000000010100111010101111100110011000111011011010100011001001011011000111101000011000010001011111110010100001001011101110001000001000011101000011110010000;
XPCT = 108'b001101110100000100001110100011110010110011111000100100011111111100011011000110110110111011111111010110111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27200

pattern = 136; // 27200
ALLPIS = 207'b010101000011011000001110010010001100110100010011011100010101001000110000000001100011110000000010110010100100100001100001001010000110000000110111011010110111110001011011100101101101101000010100101000111101101;
XPCT = 108'b001100101110110100001010010100111101110011111001111110001111011110101111010110000001110000011111110000101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27400

pattern = 137; // 27400
ALLPIS = 207'b001111011100000110110001001111100001011100101100001100011100111100001100000010100000001010101011101000110001111000010011100011010011000100000001111010101100011000010101000110010000000001001110010110011011110;
XPCT = 108'b000000110000000000100111001010011011011101111001011010000000110001111100000011111111101111000000000101011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27600

pattern = 138; // 27600
ALLPIS = 207'b110111010010011000100010010110000100011100010110101001000001000000000111101010100101000100111111011010101010000001001010001111100100111001100101011110100111100000001000011000111010010111111101111000100100100;
XPCT = 108'b110011001101001011111110111100100100001011111111011011000000000111111110011000001000100000111111001001111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27800

pattern = 139; // 27800
ALLPIS = 207'b010101000110110101101001111111111011000110100000001111010100100001111010101111001100101111010011000010110010110001010010101001011111100110000001100100010001101101100011001000011110000111010010010001001001001;
XPCT = 108'b001001000111000011101001001001001001111011111011111110010000101011011110100001001110100100111110001110100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28000

pattern = 140; // 28000
ALLPIS = 207'b100001100110010010100101111110101010011010111001110010111001000111101101000000100100011010101011100011011010011101100101011101001111011001111001110010101001101011010100100100000010110011011101000000100110001;
XPCT = 108'b110100100001011001101110100000100110100001110101111111111111110000111111011100000101111111100001110000010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28200

pattern = 141; // 28200
ALLPIS = 207'b110101010101000001100011000101010001110001011101010010010011110001101101111101001010011101111001101010110101001101000110100000011010011110100000101001110010001100111100000110011101001101001100011011100011101;
XPCT = 108'b110000110110100110100110001111100011101010111101111111101111000000001101110111101001110111011110010011000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28400

pattern = 142; // 28400
ALLPIS = 207'b011110001000110100000111001111011100111100010010100011101000011000111111110100110010001000101111000111111100001110110100011000001000010001011101100100101000000000111101011110101101000100000100111101110100001;
XPCT = 108'b000011111110100010000010011101110100010111111011011010000000000101001010101011000001100111111110101100110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28600

pattern = 143; // 28600
ALLPIS = 207'b100010011111001111000110011000001010100000110000010011100101011101110010001011000110001011001000000010100001011011011011101110101000101001011101100011010100101101111000101100111001010100100110101110010100101;
XPCT = 108'b110101101100101010010011010110010100001101111110000001101111001000001111111111100100110100011110101010101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28800

pattern = 144; // 28800
ALLPIS = 207'b000011000111111000001010000000101101000100110011101111110101001010110110110100010101111010010100100110000001010001100111010010010111000011000010100011111100100110100111000000110010001010100000111000011000111;
XPCT = 108'b001000001001000101010000011100011000011011111011010000001111010101101111101100001001111101111111010100011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29000

pattern = 145; // 29000
ALLPIS = 207'b111000110100101000010111111001101000101011111011100110000001000101111000100010001010000101010000100111110010111100001011010000110101000101010100111001011011000010111001010000110011111111001100100101101111110;
XPCT = 108'b110010001001111111100110010001101111111111111101111111001001001010010100111111111010111111100000001101100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29200

pattern = 146; // 29200
ALLPIS = 207'b001000100000011101000001010010100111001001101111001100000100011111111001011100111111001010011111110100010011001000110101011001110111011001010001100110100101000101011101011010011101001101101001110010001000001;
XPCT = 108'b000011010110100110110100111010001000111001111000100100001111111000001111100100100011110011100001100001111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29400

pattern = 147; // 29400
ALLPIS = 207'b011001010100111110110101011101000010011101000110011111001101111100100100001110011011010011111100100000000110010101001111010000110000101011000011101111010000100111010011111001101111000111000111111000001010001;
XPCT = 108'b001111001111100011100011111100001010110011111011111110010000111000101110100011001101100000111111110100100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29600

pattern = 148; // 29600
ALLPIS = 207'b011001100100000111001110000011100001100010010001011110100011000110110110011111101011001111000111100011111111010110100001000111100000101001100011100101001001011110001111101001100100111111011100000110000101001;
XPCT = 108'b001101001010011111101110000010000101110111111001111110010000111101001110110010011100101111111110011010000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29800

pattern = 149; // 29800
ALLPIS = 207'b001011010010101010010011101110010101010001110100000110001001111000101010001011001010000000000000101110000001001110100010110101101001110110011110000000110010011100100001000100101001011000110000001011101011101;
XPCT = 108'b000000101100101100011000000111101011010001111001011010001111100110011111000100011001110110100001001101001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30000

pattern = 150; // 30000
ALLPIS = 207'b011010010100001111101100001011011011001001001110111110110110011011000000101011111111110011000001101111111100011111011010101110101010011100011000010100111001111100110011000000000001001000001001100101000001010;
XPCT = 108'b001000000000100100000100110001000001010111110001011010011001010101011110101100001111111011000001101011011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30200

pattern = 151; // 30200
ALLPIS = 207'b010111001000001111101110100110001101010010111000010110101111110001001000010010100001001010000110101000010101101010110111100010110000110001010010111100000011001100010011000101011000000111101011010011011101001;
XPCT = 108'b001000100100000011110101101011011101011011111001011010011111011000011111100111110101110001000000001000011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30400

pattern = 152; // 30400
ALLPIS = 207'b100101000000000101000001100001101111100110110011101010101111110100111111001110101010011001101011110101110011010100010011111100110011100100011000111000110100011111011001111001001011111111111110000101001111001;
XPCT = 108'b110111000101111111111111000001001111110101110100100101110000111111110110010011010011101010111110101010000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30600

pattern = 153; // 30600
ALLPIS = 207'b010100110110110010011111100000001000010000011000110110000000011110011100100110011111001000011000001101111011101111011000110010011010010111101100010011100110111100111111011111000011110011101110111100110111000;
XPCT = 108'b001011110001111001110111011100110111110111011001111110011111000000011111000100010011111100000001010010001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30800

pattern = 154; // 30800
ALLPIS = 207'b000101100000110101101111011011100001110001110110001100110010011110110001100100111000101011001101001100110001010011000010110110001111010010010011011100001001100110010001101111110000000000100101101010111110101;
XPCT = 108'b000101111000000000010010110110111110111011111001110100000110110111111111111001111111100011111111110010110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31000

pattern = 155; // 31000
ALLPIS = 207'b110011101111101011111100010011000110010001010000010011011011001101101000111011010001100110001001100100010111110001101000101001101100011010110010100011111001100101010000110000110001111010011101011100010110010;
XPCT = 108'b110110001000111101001110101100010110001110101111011011011001011010111110000110010100110101011111010001110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31200

pattern = 156; // 31200
ALLPIS = 207'b010111110011000110011001110110000010110110001110110000001000001101110001001101000111101110001010000001011011011101001110111110100000000010011010011001100101011100110011110101101100011101101101001110011001010;
XPCT = 108'b001110101110001110110110100110011001010111111001011010011111111000101111100101000011110110011000000000010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31400

pattern = 157; // 31400
ALLPIS = 207'b011010001100111010100010010011010011001000011101010101110010101100101000011110010101001100001101011111100011110110011011100110011001010100010101101101110111001111001111111100000011111101101010101101000011101;
XPCT = 108'b001111100001111110110101010101000011010111011011011010000110110001101111111011111111101111111111011111000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31600

pattern = 158; // 31600
ALLPIS = 207'b111011110101101111001111011100100110100001001111111111000011011110101101011101101110101000111100010010101110010100000010001101001100011001000000111011010011101011110001110010011010001011100000111000100101010;
XPCT = 108'b110110010101000101110000011100100101011011111111011011111111100100101111110110001100110010000000111100100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31800

pattern = 159; // 31800
ALLPIS = 207'b110010111001100000000101100101000001101111010010111101110100000000011100000100010001111000000010000011110100000101110101001111100000010101000000000001001110011000100100010101000110101101010010100111011000011;
XPCT = 108'b110010100011010110101001010011011000000111111111011011111111010000110101010101111001110010111000111011011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32000

pattern = 160; // 32000
ALLPIS = 207'b110011000011111010010000000000010111010101111110000010010010100000100000010010011111100010111110100001111001100010101010101000011111100110000101111111000100001011110011010111100101001000100001010001010101100;
XPCT = 108'b111010111010100100010000101001010101010011111101011011001111101001101111100101000100110101111110100110110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32200

pattern = 161; // 32200
ALLPIS = 207'b101011011001101001100010111100001110000111011010100011011110100011011000011101001100000000111001010101010101000011100001111010010011100010010010101001101001000011101101111010011000100011111111111010010101000;
XPCT = 108'b110111010100010001111111111110010101011001111110001011011111001101001111101110101010110011111001111111100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32400

pattern = 162; // 32400
ALLPIS = 207'b101001110100011110010110011100001110000110000001010101011011001111010010011101000100110111011110001110000111011101001100000010111010011000100011001101001100111100101001101111101101001010001100110001100101101;
XPCT = 108'b110101111110100101000110011001100101110001111110101111000000000001111110100010010110101111111110110001001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32600

pattern = 163; // 32600
ALLPIS = 207'b111110100101111111010000010100100010111010000010010101000100100010100010001000011001111001011100001101101011111000011000111110000100001011100001110101111100010010111001000101110000000101011011001000110010001;
XPCT = 108'b110000101000000010101101100100110010011011111111011011111111110101100001101111111101110111011001110000111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32800

pattern = 164; // 32800
ALLPIS = 207'b010101000000100001001111001010001011010111000010010110000001101110101111100011000100010010001000110000010001110101011101111001001011111011100011100110010100111000001101100011100100110100110010101101101010111;
XPCT = 108'b000100011010011010011001010101101010110111111001111110000110010111100111001000101101100001011001111100011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33000

pattern = 165; // 33000
ALLPIS = 207'b001000100100010001000110110010010101101110100011001111000000100100000011001100101111100101001101100000001111000101101111110010000100101101010001000110011001001010100110111111010011101000101011101111000111100;
XPCT = 108'b001111110001110100010101110111000111101101111011111110001111011101010101010111010000111001100001101001100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33200

pattern = 166; // 33200
ALLPIS = 207'b101100000100111010010000011010100110100100001111111110111110011100101000010101101100110100000111100100011011100001111000001000011110010111110100010100110010101011111100100111010100001100011000100010100110000;
XPCT = 108'b110100110010000110001100010010100110101000111100101111000000001010001110010000011110100100111111010110011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33400

pattern = 167; // 33400
ALLPIS = 207'b010001000100110010110111000011011001000100111101110010000001011100010001101111110000011101000011110100010100101101000110000101100100001100111100010001111111111010000101001000010100001111101111101011101000001;
XPCT = 108'b000001000010000111110111110111101000111011111001111110010110110001111111111011011010100010111111010111100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33600

pattern = 168; // 33600
ALLPIS = 207'b000110111011011100001001111011010101100110101010011100010010100010001111100111100001110000001111001110110110110100101111111111100110110011000101111101001101110110111000111101111010001000010100100100001001101;
XPCT = 108'b000111101101000100001010010000001001001111000000001010001111110101011111011110100010111011111111010010001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33800

pattern = 169; // 33800
ALLPIS = 207'b111011001110001100111111010000111000110111101110001101111111111000111100110100000011111011110010000100000100100001001101110000001101000010110111010111111111000101011011101101110010011101100010110011101011011;
XPCT = 108'b111101101001001110110001011011101011011011111111011011110000001111110110000011101111100001111001111111110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34000

pattern = 170; // 34000
ALLPIS = 207'b100001011100011100010111001111011010001110101101001111111110001010110011101111100000101111011100011101110101011001011000000000010101111001101100011001011010101011000101101111010110111010000001110110010100110;
XPCT = 108'b110101110011011101000000111010010100111101111111110101100110101111001111101010011011100110100001111111000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34200

pattern = 171; // 34200
ALLPIS = 207'b110011011011101100000011101000000010111010110000100101100010011101010001000001100110000011100110111111101000010111111111001001101011111110000010010110011000110110101000111010010011000100110100101011111111001;
XPCT = 108'b110111010001100010011010010111111111001011111111011011011111101011101111000110011001111101111000110100100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34400

pattern = 172; // 34400
ALLPIS = 207'b001111001111011110000010011000101110000100111011010101101000101010100110011110011110011010001110001111101000000100100100100011111110110010110100011011010101100101110001101111001100100001001010010000100100101;
XPCT = 108'b000101110110010000100101001000100100010001011011011010001111000111011111000100110100111111111000110111111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34600

pattern = 173; // 34600
ALLPIS = 207'b111000000100101000100100111010001010011001110100010001100101011101111100000000100111000001010011100011101100100100001110101111001010100101101000111011000000110111000110010010010011001100111001100001001001101;
XPCT = 108'b111010010001100110011100110001001001101011111111111111011111100111100001010100001001110011000001100100110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34800

pattern = 174; // 34800
ALLPIS = 207'b100011110100111010000001100110111111111111101000001101011111110111010100011001110000101100011100011010110010101011100111101011100110100110000001111101111001000101100001100110000010111011001110111110011010001;
XPCT = 108'b110100110001011101100111011110011010010101111111011011111001100001100110111111000100111111000000011001001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35000

      $display("// %t : Simulation of %0d patterns completed with %0d errors\n", $time, pattern+1, nofails);
      if (verbose >=2) $finish(2);
      /* else */ $finish(0);
   end
endmodule
