// Verilog pattern output written by  TetraMAX (TM)  B-2008.09-SP2-i081128_181834 
// Date: Wed Jul  6 12:09:28 2011
// Module tested: c7552

//     Uncollapsed Stuck Fault Summary Report
// -----------------------------------------------
// fault class                     code   #faults
// ------------------------------  ----  ---------
// Detected                         DT       6450
// Possibly detected                PT          0
// Undetectable                     UD          0
// ATPG untestable                  AU          0
// Not detected                     ND        438
// -----------------------------------------------
// total faults                              6888
// test coverage                            93.64%
// -----------------------------------------------
// 
//            Pattern Summary Report
// -----------------------------------------------
// #internal patterns                         148
//     #basic_scan patterns                   148
// -----------------------------------------------
// 
// There are no rule fails
// There are no clocks
// There are no constraint ports
// There are no equivalent pins
// There are no net connections

`timescale 1 ns / 1 ns

//
// --- NOTE: Remove the comment to define 'tmax_iddq' to activate processing of IDDQ events
//     Or use '+define+tmax_iddq' on the verilog compile line
//
//`define tmax_iddq

module AAA_tmax_testbench_1_16 ;
   parameter NAMELENGTH = 200; // max length of names reported in fails
   integer nofails, bit, pattern, lastpattern;
   integer error_banner; // flag for tracking displayed error banner
   integer loads;        // number of load_unloads for current pattern
   integer patm1;        // pattern - 1
   integer patp1;        // pattern + lastpattern
   integer prev_pat;     // previous pattern number
   integer report_interval; // report pattern progress every Nth pattern
   integer verbose;      // message verbosity level
   parameter NINPUTS = 207, NOUTPUTS = 108;
   wire [0:NOUTPUTS-1] PO; reg [0:NOUTPUTS-1] ALLPOS, XPCT, MASK;
   reg [0:NINPUTS-1] PI, ALLPIS;
   reg [0:8*(NAMELENGTH-1)] POnames [0:NOUTPUTS-1];
   event IDDQ;

   wire N1;
   wire N5;
   wire N9;
   wire N12;
   wire N15;
   wire N18;
   wire N23;
   wire N26;
   wire N29;
   wire N32;
   wire N35;
   wire N38;
   wire N41;
   wire N44;
   wire N47;
   wire N50;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N69;
   wire N70;
   wire N73;
   wire N74;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N82;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N94;
   wire N97;
   wire N100;
   wire N103;
   wire N106;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N118;
   wire N121;
   wire N124;
   wire N127;
   wire N130;
   wire N133;
   wire N134;
   wire N135;
   wire N138;
   wire N141;
   wire N144;
   wire N147;
   wire N150;
   wire N151;
   wire N152;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N178;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire N185;
   wire N186;
   wire N187;
   wire N188;
   wire N189;
   wire N190;
   wire N191;
   wire N192;
   wire N193;
   wire N194;
   wire N195;
   wire N196;
   wire N197;
   wire N198;
   wire N199;
   wire N200;
   wire N201;
   wire N202;
   wire N203;
   wire N204;
   wire N205;
   wire N206;
   wire N207;
   wire N208;
   wire N209;
   wire N210;
   wire N211;
   wire N212;
   wire N213;
   wire N214;
   wire N215;
   wire N216;
   wire N217;
   wire N218;
   wire N219;
   wire N220;
   wire N221;
   wire N222;
   wire N223;
   wire N224;
   wire N225;
   wire N226;
   wire N227;
   wire N228;
   wire N229;
   wire N230;
   wire N231;
   wire N232;
   wire N233;
   wire N234;
   wire N235;
   wire N236;
   wire N237;
   wire N238;
   wire N239;
   wire N240;
   wire N242;
   wire N245;
   wire N248;
   wire N251;
   wire N254;
   wire N257;
   wire N260;
   wire N263;
   wire N267;
   wire N271;
   wire N274;
   wire N277;
   wire N280;
   wire N283;
   wire N286;
   wire N289;
   wire N293;
   wire N296;
   wire N299;
   wire N303;
   wire N307;
   wire N310;
   wire N313;
   wire N316;
   wire N319;
   wire N322;
   wire N325;
   wire N328;
   wire N331;
   wire N334;
   wire N337;
   wire N340;
   wire N343;
   wire N346;
   wire N349;
   wire N352;
   wire N355;
   wire N358;
   wire N361;
   wire N364;
   wire N367;
   wire N382;
   wire N241_I;
   wire N387;
   wire N388;
   wire N478;
   wire N482;
   wire N484;
   wire N486;
   wire N489;
   wire N492;
   wire N501;
   wire N505;
   wire N507;
   wire N509;
   wire N511;
   wire N513;
   wire N515;
   wire N517;
   wire N519;
   wire N535;
   wire N537;
   wire N539;
   wire N541;
   wire N543;
   wire N545;
   wire N547;
   wire N549;
   wire N551;
   wire N553;
   wire N556;
   wire N559;
   wire N561;
   wire N563;
   wire N565;
   wire N567;
   wire N569;
   wire N571;
   wire N573;
   wire N582;
   wire N643;
   wire N707;
   wire N813;
   wire N881;
   wire N882;
   wire N883;
   wire N884;
   wire N885;
   wire N889;
   wire N945;
   wire N1110;
   wire N1111;
   wire N1112;
   wire N1113;
   wire N1114;
   wire N1489;
   wire N1490;
   wire N1781;
   wire N10025;
   wire N10101;
   wire N10102;
   wire N10103;
   wire N10104;
   wire N10109;
   wire N10110;
   wire N10111;
   wire N10112;
   wire N10350;
   wire N10351;
   wire N10352;
   wire N10353;
   wire N10574;
   wire N10575;
   wire N10576;
   wire N10628;
   wire N10632;
   wire N10641;
   wire N10704;
   wire N10706;
   wire N10711;
   wire N10712;
   wire N10713;
   wire N10714;
   wire N10715;
   wire N10716;
   wire N10717;
   wire N10718;
   wire N10729;
   wire N10759;
   wire N10760;
   wire N10761;
   wire N10762;
   wire N10763;
   wire N10827;
   wire N10837;
   wire N10838;
   wire N10839;
   wire N10840;
   wire N10868;
   wire N10869;
   wire N10870;
   wire N10871;
   wire N10905;
   wire N10906;
   wire N10907;
   wire N10908;
   wire N11333;
   wire N11334;
   wire N11340;
   wire N11342;
   wire N241_O;

   // map PI[] vector to DUT inputs and bidis
   assign N1 = PI[0];
   assign N5 = PI[1];
   assign N9 = PI[2];
   assign N12 = PI[3];
   assign N15 = PI[4];
   assign N18 = PI[5];
   assign N23 = PI[6];
   assign N26 = PI[7];
   assign N29 = PI[8];
   assign N32 = PI[9];
   assign N35 = PI[10];
   assign N38 = PI[11];
   assign N41 = PI[12];
   assign N44 = PI[13];
   assign N47 = PI[14];
   assign N50 = PI[15];
   assign N53 = PI[16];
   assign N54 = PI[17];
   assign N55 = PI[18];
   assign N56 = PI[19];
   assign N57 = PI[20];
   assign N58 = PI[21];
   assign N59 = PI[22];
   assign N60 = PI[23];
   assign N61 = PI[24];
   assign N62 = PI[25];
   assign N63 = PI[26];
   assign N64 = PI[27];
   assign N65 = PI[28];
   assign N66 = PI[29];
   assign N69 = PI[30];
   assign N70 = PI[31];
   assign N73 = PI[32];
   assign N74 = PI[33];
   assign N75 = PI[34];
   assign N76 = PI[35];
   assign N77 = PI[36];
   assign N78 = PI[37];
   assign N79 = PI[38];
   assign N80 = PI[39];
   assign N81 = PI[40];
   assign N82 = PI[41];
   assign N83 = PI[42];
   assign N84 = PI[43];
   assign N85 = PI[44];
   assign N86 = PI[45];
   assign N87 = PI[46];
   assign N88 = PI[47];
   assign N89 = PI[48];
   assign N94 = PI[49];
   assign N97 = PI[50];
   assign N100 = PI[51];
   assign N103 = PI[52];
   assign N106 = PI[53];
   assign N109 = PI[54];
   assign N110 = PI[55];
   assign N111 = PI[56];
   assign N112 = PI[57];
   assign N113 = PI[58];
   assign N114 = PI[59];
   assign N115 = PI[60];
   assign N118 = PI[61];
   assign N121 = PI[62];
   assign N124 = PI[63];
   assign N127 = PI[64];
   assign N130 = PI[65];
   assign N133 = PI[66];
   assign N134 = PI[67];
   assign N135 = PI[68];
   assign N138 = PI[69];
   assign N141 = PI[70];
   assign N144 = PI[71];
   assign N147 = PI[72];
   assign N150 = PI[73];
   assign N151 = PI[74];
   assign N152 = PI[75];
   assign N153 = PI[76];
   assign N154 = PI[77];
   assign N155 = PI[78];
   assign N156 = PI[79];
   assign N157 = PI[80];
   assign N158 = PI[81];
   assign N159 = PI[82];
   assign N160 = PI[83];
   assign N161 = PI[84];
   assign N162 = PI[85];
   assign N163 = PI[86];
   assign N164 = PI[87];
   assign N165 = PI[88];
   assign N166 = PI[89];
   assign N167 = PI[90];
   assign N168 = PI[91];
   assign N169 = PI[92];
   assign N170 = PI[93];
   assign N171 = PI[94];
   assign N172 = PI[95];
   assign N173 = PI[96];
   assign N174 = PI[97];
   assign N175 = PI[98];
   assign N176 = PI[99];
   assign N177 = PI[100];
   assign N178 = PI[101];
   assign N179 = PI[102];
   assign N180 = PI[103];
   assign N181 = PI[104];
   assign N182 = PI[105];
   assign N183 = PI[106];
   assign N184 = PI[107];
   assign N185 = PI[108];
   assign N186 = PI[109];
   assign N187 = PI[110];
   assign N188 = PI[111];
   assign N189 = PI[112];
   assign N190 = PI[113];
   assign N191 = PI[114];
   assign N192 = PI[115];
   assign N193 = PI[116];
   assign N194 = PI[117];
   assign N195 = PI[118];
   assign N196 = PI[119];
   assign N197 = PI[120];
   assign N198 = PI[121];
   assign N199 = PI[122];
   assign N200 = PI[123];
   assign N201 = PI[124];
   assign N202 = PI[125];
   assign N203 = PI[126];
   assign N204 = PI[127];
   assign N205 = PI[128];
   assign N206 = PI[129];
   assign N207 = PI[130];
   assign N208 = PI[131];
   assign N209 = PI[132];
   assign N210 = PI[133];
   assign N211 = PI[134];
   assign N212 = PI[135];
   assign N213 = PI[136];
   assign N214 = PI[137];
   assign N215 = PI[138];
   assign N216 = PI[139];
   assign N217 = PI[140];
   assign N218 = PI[141];
   assign N219 = PI[142];
   assign N220 = PI[143];
   assign N221 = PI[144];
   assign N222 = PI[145];
   assign N223 = PI[146];
   assign N224 = PI[147];
   assign N225 = PI[148];
   assign N226 = PI[149];
   assign N227 = PI[150];
   assign N228 = PI[151];
   assign N229 = PI[152];
   assign N230 = PI[153];
   assign N231 = PI[154];
   assign N232 = PI[155];
   assign N233 = PI[156];
   assign N234 = PI[157];
   assign N235 = PI[158];
   assign N236 = PI[159];
   assign N237 = PI[160];
   assign N238 = PI[161];
   assign N239 = PI[162];
   assign N240 = PI[163];
   assign N242 = PI[164];
   assign N245 = PI[165];
   assign N248 = PI[166];
   assign N251 = PI[167];
   assign N254 = PI[168];
   assign N257 = PI[169];
   assign N260 = PI[170];
   assign N263 = PI[171];
   assign N267 = PI[172];
   assign N271 = PI[173];
   assign N274 = PI[174];
   assign N277 = PI[175];
   assign N280 = PI[176];
   assign N283 = PI[177];
   assign N286 = PI[178];
   assign N289 = PI[179];
   assign N293 = PI[180];
   assign N296 = PI[181];
   assign N299 = PI[182];
   assign N303 = PI[183];
   assign N307 = PI[184];
   assign N310 = PI[185];
   assign N313 = PI[186];
   assign N316 = PI[187];
   assign N319 = PI[188];
   assign N322 = PI[189];
   assign N325 = PI[190];
   assign N328 = PI[191];
   assign N331 = PI[192];
   assign N334 = PI[193];
   assign N337 = PI[194];
   assign N340 = PI[195];
   assign N343 = PI[196];
   assign N346 = PI[197];
   assign N349 = PI[198];
   assign N352 = PI[199];
   assign N355 = PI[200];
   assign N358 = PI[201];
   assign N361 = PI[202];
   assign N364 = PI[203];
   assign N367 = PI[204];
   assign N382 = PI[205];
   assign N241_I = PI[206];

   // map DUT outputs and bidis to PO[] vector
   assign
      PO[0] = N387 ,
      PO[1] = N388 ,
      PO[2] = N478 ,
      PO[3] = N482 ,
      PO[4] = N484 ,
      PO[5] = N486 ,
      PO[6] = N489 ,
      PO[7] = N492 ,
      PO[8] = N501 ,
      PO[9] = N505 ,
      PO[10] = N507 ,
      PO[11] = N509 ,
      PO[12] = N511 ,
      PO[13] = N513 ,
      PO[14] = N515 ,
      PO[15] = N517 ,
      PO[16] = N519 ,
      PO[17] = N535 ,
      PO[18] = N537 ,
      PO[19] = N539 ,
      PO[20] = N541 ,
      PO[21] = N543 ,
      PO[22] = N545 ,
      PO[23] = N547 ,
      PO[24] = N549 ,
      PO[25] = N551 ,
      PO[26] = N553 ,
      PO[27] = N556 ,
      PO[28] = N559 ,
      PO[29] = N561 ,
      PO[30] = N563 ,
      PO[31] = N565 ;
   assign
      PO[32] = N567 ,
      PO[33] = N569 ,
      PO[34] = N571 ,
      PO[35] = N573 ,
      PO[36] = N582 ,
      PO[37] = N643 ,
      PO[38] = N707 ,
      PO[39] = N813 ,
      PO[40] = N881 ,
      PO[41] = N882 ,
      PO[42] = N883 ,
      PO[43] = N884 ,
      PO[44] = N885 ,
      PO[45] = N889 ,
      PO[46] = N945 ,
      PO[47] = N1110 ,
      PO[48] = N1111 ,
      PO[49] = N1112 ,
      PO[50] = N1113 ,
      PO[51] = N1114 ,
      PO[52] = N1489 ,
      PO[53] = N1490 ,
      PO[54] = N1781 ,
      PO[55] = N10025 ,
      PO[56] = N10101 ,
      PO[57] = N10102 ,
      PO[58] = N10103 ,
      PO[59] = N10104 ,
      PO[60] = N10109 ,
      PO[61] = N10110 ,
      PO[62] = N10111 ,
      PO[63] = N10112 ;
   assign
      PO[64] = N10350 ,
      PO[65] = N10351 ,
      PO[66] = N10352 ,
      PO[67] = N10353 ,
      PO[68] = N10574 ,
      PO[69] = N10575 ,
      PO[70] = N10576 ,
      PO[71] = N10628 ,
      PO[72] = N10632 ,
      PO[73] = N10641 ,
      PO[74] = N10704 ,
      PO[75] = N10706 ,
      PO[76] = N10711 ,
      PO[77] = N10712 ,
      PO[78] = N10713 ,
      PO[79] = N10714 ,
      PO[80] = N10715 ,
      PO[81] = N10716 ,
      PO[82] = N10717 ,
      PO[83] = N10718 ,
      PO[84] = N10729 ,
      PO[85] = N10759 ,
      PO[86] = N10760 ,
      PO[87] = N10761 ,
      PO[88] = N10762 ,
      PO[89] = N10763 ,
      PO[90] = N10827 ,
      PO[91] = N10837 ,
      PO[92] = N10838 ,
      PO[93] = N10839 ,
      PO[94] = N10840 ,
      PO[95] = N10868 ;
   assign
      PO[96] = N10869 ,
      PO[97] = N10870 ,
      PO[98] = N10871 ,
      PO[99] = N10905 ,
      PO[100] = N10906 ,
      PO[101] = N10907 ,
      PO[102] = N10908 ,
      PO[103] = N11333 ,
      PO[104] = N11334 ,
      PO[105] = N11340 ,
      PO[106] = N11342 ,
      PO[107] = N241_O ;

   // instantiate the design into the testbench
   c7552 dut (
      .N1(N1),
      .N5(N5),
      .N9(N9),
      .N12(N12),
      .N15(N15),
      .N18(N18),
      .N23(N23),
      .N26(N26),
      .N29(N29),
      .N32(N32),
      .N35(N35),
      .N38(N38),
      .N41(N41),
      .N44(N44),
      .N47(N47),
      .N50(N50),
      .N53(N53),
      .N54(N54),
      .N55(N55),
      .N56(N56),
      .N57(N57),
      .N58(N58),
      .N59(N59),
      .N60(N60),
      .N61(N61),
      .N62(N62),
      .N63(N63),
      .N64(N64),
      .N65(N65),
      .N66(N66),
      .N69(N69),
      .N70(N70),
      .N73(N73),
      .N74(N74),
      .N75(N75),
      .N76(N76),
      .N77(N77),
      .N78(N78),
      .N79(N79),
      .N80(N80),
      .N81(N81),
      .N82(N82),
      .N83(N83),
      .N84(N84),
      .N85(N85),
      .N86(N86),
      .N87(N87),
      .N88(N88),
      .N89(N89),
      .N94(N94),
      .N97(N97),
      .N100(N100),
      .N103(N103),
      .N106(N106),
      .N109(N109),
      .N110(N110),
      .N111(N111),
      .N112(N112),
      .N113(N113),
      .N114(N114),
      .N115(N115),
      .N118(N118),
      .N121(N121),
      .N124(N124),
      .N127(N127),
      .N130(N130),
      .N133(N133),
      .N134(N134),
      .N135(N135),
      .N138(N138),
      .N141(N141),
      .N144(N144),
      .N147(N147),
      .N150(N150),
      .N151(N151),
      .N152(N152),
      .N153(N153),
      .N154(N154),
      .N155(N155),
      .N156(N156),
      .N157(N157),
      .N158(N158),
      .N159(N159),
      .N160(N160),
      .N161(N161),
      .N162(N162),
      .N163(N163),
      .N164(N164),
      .N165(N165),
      .N166(N166),
      .N167(N167),
      .N168(N168),
      .N169(N169),
      .N170(N170),
      .N171(N171),
      .N172(N172),
      .N173(N173),
      .N174(N174),
      .N175(N175),
      .N176(N176),
      .N177(N177),
      .N178(N178),
      .N179(N179),
      .N180(N180),
      .N181(N181),
      .N182(N182),
      .N183(N183),
      .N184(N184),
      .N185(N185),
      .N186(N186),
      .N187(N187),
      .N188(N188),
      .N189(N189),
      .N190(N190),
      .N191(N191),
      .N192(N192),
      .N193(N193),
      .N194(N194),
      .N195(N195),
      .N196(N196),
      .N197(N197),
      .N198(N198),
      .N199(N199),
      .N200(N200),
      .N201(N201),
      .N202(N202),
      .N203(N203),
      .N204(N204),
      .N205(N205),
      .N206(N206),
      .N207(N207),
      .N208(N208),
      .N209(N209),
      .N210(N210),
      .N211(N211),
      .N212(N212),
      .N213(N213),
      .N214(N214),
      .N215(N215),
      .N216(N216),
      .N217(N217),
      .N218(N218),
      .N219(N219),
      .N220(N220),
      .N221(N221),
      .N222(N222),
      .N223(N223),
      .N224(N224),
      .N225(N225),
      .N226(N226),
      .N227(N227),
      .N228(N228),
      .N229(N229),
      .N230(N230),
      .N231(N231),
      .N232(N232),
      .N233(N233),
      .N234(N234),
      .N235(N235),
      .N236(N236),
      .N237(N237),
      .N238(N238),
      .N239(N239),
      .N240(N240),
      .N242(N242),
      .N245(N245),
      .N248(N248),
      .N251(N251),
      .N254(N254),
      .N257(N257),
      .N260(N260),
      .N263(N263),
      .N267(N267),
      .N271(N271),
      .N274(N274),
      .N277(N277),
      .N280(N280),
      .N283(N283),
      .N286(N286),
      .N289(N289),
      .N293(N293),
      .N296(N296),
      .N299(N299),
      .N303(N303),
      .N307(N307),
      .N310(N310),
      .N313(N313),
      .N316(N316),
      .N319(N319),
      .N322(N322),
      .N325(N325),
      .N328(N328),
      .N331(N331),
      .N334(N334),
      .N337(N337),
      .N340(N340),
      .N343(N343),
      .N346(N346),
      .N349(N349),
      .N352(N352),
      .N355(N355),
      .N358(N358),
      .N361(N361),
      .N364(N364),
      .N367(N367),
      .N382(N382),
      .N241_I(N241_I),
      .N387(N387),
      .N388(N388),
      .N478(N478),
      .N482(N482),
      .N484(N484),
      .N486(N486),
      .N489(N489),
      .N492(N492),
      .N501(N501),
      .N505(N505),
      .N507(N507),
      .N509(N509),
      .N511(N511),
      .N513(N513),
      .N515(N515),
      .N517(N517),
      .N519(N519),
      .N535(N535),
      .N537(N537),
      .N539(N539),
      .N541(N541),
      .N543(N543),
      .N545(N545),
      .N547(N547),
      .N549(N549),
      .N551(N551),
      .N553(N553),
      .N556(N556),
      .N559(N559),
      .N561(N561),
      .N563(N563),
      .N565(N565),
      .N567(N567),
      .N569(N569),
      .N571(N571),
      .N573(N573),
      .N582(N582),
      .N643(N643),
      .N707(N707),
      .N813(N813),
      .N881(N881),
      .N882(N882),
      .N883(N883),
      .N884(N884),
      .N885(N885),
      .N889(N889),
      .N945(N945),
      .N1110(N1110),
      .N1111(N1111),
      .N1112(N1112),
      .N1113(N1113),
      .N1114(N1114),
      .N1489(N1489),
      .N1490(N1490),
      .N1781(N1781),
      .N10025(N10025),
      .N10101(N10101),
      .N10102(N10102),
      .N10103(N10103),
      .N10104(N10104),
      .N10109(N10109),
      .N10110(N10110),
      .N10111(N10111),
      .N10112(N10112),
      .N10350(N10350),
      .N10351(N10351),
      .N10352(N10352),
      .N10353(N10353),
      .N10574(N10574),
      .N10575(N10575),
      .N10576(N10576),
      .N10628(N10628),
      .N10632(N10632),
      .N10641(N10641),
      .N10704(N10704),
      .N10706(N10706),
      .N10711(N10711),
      .N10712(N10712),
      .N10713(N10713),
      .N10714(N10714),
      .N10715(N10715),
      .N10716(N10716),
      .N10717(N10717),
      .N10718(N10718),
      .N10729(N10729),
      .N10759(N10759),
      .N10760(N10760),
      .N10761(N10761),
      .N10762(N10762),
      .N10763(N10763),
      .N10827(N10827),
      .N10837(N10837),
      .N10838(N10838),
      .N10839(N10839),
      .N10840(N10840),
      .N10868(N10868),
      .N10869(N10869),
      .N10870(N10870),
      .N10871(N10871),
      .N10905(N10905),
      .N10906(N10906),
      .N10907(N10907),
      .N10908(N10908),
      .N11333(N11333),
      .N11334(N11334),
      .N11340(N11340),
      .N11342(N11342),
      .N241_O(N241_O)   );


   integer errshown;
   event measurePO;
   always @ measurePO begin
      if (((XPCT&MASK) !== (ALLPOS&MASK)) || (XPCT !== (~(~XPCT)))) begin
         errshown = 0;
         for (bit = 0; bit < NOUTPUTS; bit=bit + 1) begin
            if (MASK[bit]==1'b1) begin
               if (XPCT[bit] !== ALLPOS[bit]) begin
                  if (errshown==0) $display("\n// *** ERROR during capture pattern %0d, T=%t", pattern, $time);
                  $display("  %0d %0s (exp=%b, got=%b)", pattern, POnames[bit], XPCT[bit], ALLPOS[bit]);
                  nofails = nofails + 1; errshown = 1;
               end
            end
         end
      end
   end

   event forcePI_default_WFT;
   always @ forcePI_default_WFT begin
      PI = ALLPIS;
   end
   event measurePO_default_WFT;
   always @ measurePO_default_WFT begin
      #40;
      ALLPOS = PO;
      #0; #0 -> measurePO;
      `ifdef tmax_iddq
         #0; ->IDDQ;
      `endif
   end

   always @ IDDQ begin
   `ifdef tmax_iddq
      $ssi_iddq("strobe_try");
      $ssi_iddq("status drivers leaky AAA_tmax_testbench_1_16.leaky");
   `endif
   end

   event capture;
   always @ capture begin
      ->forcePI_default_WFT;
      #100; ->measurePO_default_WFT;
   end


   initial begin

      //
      // --- establish a default time format for %t
      //
      $timeformat(-9,2," ns",18);

      //
      // --- default verbosity to 2 but also allow user override by
      //     using '+define+tmax_msg=N' on verilog compile line.
      //
      `ifdef tmax_msg
         verbose = `tmax_msg ;
      `else
         verbose = 2 ;
      `endif

      //
      // --- default pattern reporting interval to 5 but also allow user
      //     override by using '+define+tmax_rpt=N' on verilog compile line.
      //
      `ifdef tmax_rpt
         report_interval = `tmax_rpt ;
      `else
         report_interval = 5 ;
      `endif

      //
      // --- support generating Extened VCD output by using
      //     '+define+tmax_vcde' on verilog compile line.
      //
      `ifdef tmax_vcde
         // extended VCD, see IEEE Verilog P1364.1-1999 Draft 2
         if (verbose >= 2) $display("// %t : opening Extended VCD output file", $time);
         $dumpports( dut, "sim_vcde.out");
      `endif

      //
      // --- IDDQ PLI initialization
      //     User may activite by using '+define+tmax_iddq' on verilog compile line.
      //     Or by defining `tmax_iddq in this file.
      //
      `ifdef tmax_iddq
         if (verbose >= 3) $display("// %t : Initializing IDDQ PLI", $time);
         $ssi_iddq("dut AAA_tmax_testbench_1_16.dut");
         $ssi_iddq("verb on");
         $ssi_iddq("cycle 0");
         //
         // --- User may select one of the following two methods for fault seeding:
         //     #1 faults seeded by PLI (default)
         //     #2 faults supplied in a file
         //     Comment out the unused lines as needed (precede with '//').
         //     Replace the 'FAULTLIST_FILE' string with the actual file pathname.
         //
         $ssi_iddq("seed SA AAA_tmax_testbench_1_16.dut");   // no file, faults seeded by PLI
         //
         // $ssi_iddq("scope AAA_tmax_testbench_1_16.dut");   // set scope for faults from a file
         // $ssi_iddq("read_tmax FAULTLIST_FILE"); // read faults from a file
         //
      `endif

      POnames[0] = "N387";
      POnames[1] = "N388";
      POnames[2] = "N478";
      POnames[3] = "N482";
      POnames[4] = "N484";
      POnames[5] = "N486";
      POnames[6] = "N489";
      POnames[7] = "N492";
      POnames[8] = "N501";
      POnames[9] = "N505";
      POnames[10] = "N507";
      POnames[11] = "N509";
      POnames[12] = "N511";
      POnames[13] = "N513";
      POnames[14] = "N515";
      POnames[15] = "N517";
      POnames[16] = "N519";
      POnames[17] = "N535";
      POnames[18] = "N537";
      POnames[19] = "N539";
      POnames[20] = "N541";
      POnames[21] = "N543";
      POnames[22] = "N545";
      POnames[23] = "N547";
      POnames[24] = "N549";
      POnames[25] = "N551";
      POnames[26] = "N553";
      POnames[27] = "N556";
      POnames[28] = "N559";
      POnames[29] = "N561";
      POnames[30] = "N563";
      POnames[31] = "N565";
      POnames[32] = "N567";
      POnames[33] = "N569";
      POnames[34] = "N571";
      POnames[35] = "N573";
      POnames[36] = "N582";
      POnames[37] = "N643";
      POnames[38] = "N707";
      POnames[39] = "N813";
      POnames[40] = "N881";
      POnames[41] = "N882";
      POnames[42] = "N883";
      POnames[43] = "N884";
      POnames[44] = "N885";
      POnames[45] = "N889";
      POnames[46] = "N945";
      POnames[47] = "N1110";
      POnames[48] = "N1111";
      POnames[49] = "N1112";
      POnames[50] = "N1113";
      POnames[51] = "N1114";
      POnames[52] = "N1489";
      POnames[53] = "N1490";
      POnames[54] = "N1781";
      POnames[55] = "N10025";
      POnames[56] = "N10101";
      POnames[57] = "N10102";
      POnames[58] = "N10103";
      POnames[59] = "N10104";
      POnames[60] = "N10109";
      POnames[61] = "N10110";
      POnames[62] = "N10111";
      POnames[63] = "N10112";
      POnames[64] = "N10350";
      POnames[65] = "N10351";
      POnames[66] = "N10352";
      POnames[67] = "N10353";
      POnames[68] = "N10574";
      POnames[69] = "N10575";
      POnames[70] = "N10576";
      POnames[71] = "N10628";
      POnames[72] = "N10632";
      POnames[73] = "N10641";
      POnames[74] = "N10704";
      POnames[75] = "N10706";
      POnames[76] = "N10711";
      POnames[77] = "N10712";
      POnames[78] = "N10713";
      POnames[79] = "N10714";
      POnames[80] = "N10715";
      POnames[81] = "N10716";
      POnames[82] = "N10717";
      POnames[83] = "N10718";
      POnames[84] = "N10729";
      POnames[85] = "N10759";
      POnames[86] = "N10760";
      POnames[87] = "N10761";
      POnames[88] = "N10762";
      POnames[89] = "N10763";
      POnames[90] = "N10827";
      POnames[91] = "N10837";
      POnames[92] = "N10838";
      POnames[93] = "N10839";
      POnames[94] = "N10840";
      POnames[95] = "N10868";
      POnames[96] = "N10869";
      POnames[97] = "N10870";
      POnames[98] = "N10871";
      POnames[99] = "N10905";
      POnames[100] = "N10906";
      POnames[101] = "N10907";
      POnames[102] = "N10908";
      POnames[103] = "N11333";
      POnames[104] = "N11334";
      POnames[105] = "N11340";
      POnames[106] = "N11342";
      POnames[107] = "N241_O";
      nofails = 0; pattern = -1; lastpattern = 0;
      prev_pat = -2; error_banner = -2;
      /*** No test setup procedure ***/


      /*** Non-scan test ***/

      if (verbose >= 1) $display("// %t : Begin patterns, first pattern = 0", $time);
pattern = 0; // 0
ALLPIS = 207'b011100110111110010001000010000010100011111001011111101011101100010001000101001101010010011010000001111100111000101110000011010110011010111001111101000110010000011010000011101010111001100100010100100000100111;
XPCT = 108'b000011100011100110010001010000000100101111111011111110011111010101011111010101100001110011100110010000110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 200

pattern = 1; // 200
ALLPIS = 207'b001110011011111001000100001000001010001111100101111110101110110001000100010100110101001001101000000111110011100010111000001101011001101011100111110100011001000001101000001110101011100110010001010010000010011;
XPCT = 108'b000001111101110011001000101010000010000001111000001010000000100111111110110000110111100110011111010110101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 400

pattern = 2; // 400
ALLPIS = 207'b111011111010001110101010010100010001011000111001000010001010111010101010100011110000110111100100001100011110110100101100011100011111100010111100010010111110100011100100011010000010111111101010001101000101110;
XPCT = 108'b110011010001011111110101000101000101000111101101011011000000111010001010100010111111101111000110000011110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 600

pattern = 3; // 600
ALLPIS = 207'b100001001010110101011101011010011100110011010111011100011000111111011101111000010010001000100010001001101000011111100110010100111100100110010001100001101101010010100010010000010110010011010111100010100110000;
XPCT = 108'b111010000011001001101011110010100110101011111101111111111111011111011111101110110101111110100001011111101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 800

pattern = 4; // 800
ALLPIS = 207'b001100010010101000100110111101011010000110100000010011010001111101100110010101100011010111000001001011010011001010000011010000101101000100000111011000000100101010000001010101011100000101001001010101010111111;
XPCT = 108'b000010100110000010100100101001010111111101111011111110000000011010111110001011011001100111111000011101110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1000

pattern = 5; // 1000
ALLPIS = 207'b100110001001010100010011011110101101000011010000001001101000111110110011001010110001101011100000100101101001100101000001101000010110100010000011101100000010010101000000101010101110000010100100101010101011111;
XPCT = 108'b110101011111000001010010010110101011000001111111010001101111100000011111110100100100111111100110000011110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1200

pattern = 6; // 1200
ALLPIS = 207'b001111110011011000000001111111000010111110100011111001101001111101010001001100110010100110100000011101010011110111010000101110111000000110001110011110110011001001110000001000000000001101110000110001010001000;
XPCT = 108'b000001000000000110111000011001010001000001111011011010011111010100000111111100100101110100111000100000101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1400

pattern = 7; // 1400
ALLPIS = 207'b000111111001101100000000111111100001011111010001111100110100111110101000100110011001010011010000001110101001111011101000010111011100000011000111001111011001100100111000000100000000000110111000011000101000100;
XPCT = 108'b000000100000000011011100001100101000000001111000001010001111110111011001001110011100110001111111010101101110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1600

pattern = 8; // 1600
ALLPIS = 207'b111111001011000100001000001111100100110000100011000011000111111101011100111010100110111010111000001000110011111000000100010001011101010110101100001111011110110001001100011111010111001111111110101000010000101;
XPCT = 108'b110011110011100111111111010100010000001011111111011011101111001001011111010110000001110011111000111000000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1800

pattern = 9; // 1800
ALLPIS = 207'b011111100101100010000100000111110010011000010001100001100011111110101110011101010011011101011100000100011001111100000010001000101110101011010110000111101111011000100110001111101011100111111111010100001000010;
XPCT = 108'b001001111101110011111111101000001000000111111011011010010110100000011111110001100101100110111110110011100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2000

pattern = 10; // 2000
ALLPIS = 207'b101111110010110001000010000011111001001100001000110000110001111111010111001110101001101110101110000010001100111110000001000100010111010101101011000011110111101100010011000111110101110011111111101010000100001;
XPCT = 108'b111000111010111001111111110110000100011001111101011011110000110001101110001001111111101100111110010101001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2200

pattern = 11; // 2200
ALLPIS = 207'b001011001110101010101001010001101000111001001111100101000101011101100011001110111110100100000111001110100001011010110000111000111000111101111010001001001001110101011001111110101101110101011101010001000110111;
XPCT = 108'b000111111110111010101110101001000110010011111010001010000000011111001110101000111000100000000000111001000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2400

pattern = 12; // 2400
ALLPIS = 207'b011001010000100111011100111000100000000011101100001111111111001100111001001110110101000001010011101000110111101000101000000110101111001001110010101100010110111001111100100010000001110110001100001100100111100;
XPCT = 108'b000100010000111011000110000100100111100111111011111110001111110110101111010111010011111111100000111110000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2600

pattern = 13; // 2600
ALLPIS = 207'b001100101000010011101110011100010000000001110110000111111111100110011100100111011010100000101001110100011011110100010100000011010111100100111001010110001011011100111110010001000000111011000110000110010011110;
XPCT = 108'b001010000000011101100011000010010011100111111010101110010000010011010100010001011001101001111110110001110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2800

pattern = 14; // 2800
ALLPIS = 207'b111010100011111011111111011110011100011111110000111110100010010001000110111010000111000011000100110101101010111111111010011011011000100101010011000011110111101101001111010101110111010001000001100111001101000;
XPCT = 108'b111010101011101000100000110011001101011111111101011011011111101100111111100110101011111100011111000011000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3000

pattern = 15; // 3000
ALLPIS = 207'b011101010001111101111111101111001110001111111000011111010001001000100011011101000011100001100010011010110101011111111101001101101100010010101001100001111011110110100111101010111011101000100000110011100110100;
XPCT = 108'b001101011101110100010000011011100110111011111011111110001111010100111111101101010100111010111001010111101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3200

pattern = 16; // 3200
ALLPIS = 207'b010010011111001100110111100111110011011000110111110010110101000110011001000111001011100011100001000010111101101010001110111100000101011110011011011000001111111000000011101000001010111000110010111101110111101;
XPCT = 108'b001101000101011100011001011101110111010111111001011010001111100010011111001110010110111000011111011000001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3400

pattern = 17; // 3400
ALLPIS = 207'b010101111000010100010011100011101101110011010000000100000111000001000100001010001111100010100000101110111001110000110111000100110001111000000010000100110101111111010001101001010010010000111011111010111111001;
XPCT = 108'b000101000001001000011101111110111111111011111001111110010000011110001110100010100111100110111110110100000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3600

pattern = 18; // 3600
ALLPIS = 207'b001010111100001010001001110001110110111001101000000010000011100000100010000101000111110001010000010111011100111000011011100010011000111100000001000010011010111111101000110100101001001000011101111101011111100;
XPCT = 108'b000110101100100100001110111101011111000111111000001010001111000100101111111111101010111010000001101101010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3800

pattern = 19; // 3800
ALLPIS = 207'b000101011110000101000100111000111011011100110100000001000001110000010001000010100011111000101000001011101110011100001101110001001100011110000000100001001101011111110100011010010100100100001110111110101111110;
XPCT = 108'b000011010010010010000111011110101111101101111011111110000000001110001110000000001010100001000111011001000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4000

pattern = 20; // 4000
ALLPIS = 207'b000010101111000010100010011100011101101110011010000000100000111000001000100001010001111100010100000101110111001110000110111000100110001111000000010000100110101111111010001101001010010010000111011111010111111;
XPCT = 108'b001001100101001001000011101111010111000101111000001010001111110101001111010101110111111101111001000010010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4200

pattern = 21; // 4200
ALLPIS = 207'b100001010111100001010001001110001110110111001101000000010000011100000100010000101000111110001010000010111011100111000011011100010011000111100000001000010011010111111101000110100101001001000011101111101011111;
XPCT = 108'b110000111010100100100001110111101011110100111100101111101111011101101111100111011101111101100000000001100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4400

pattern = 22; // 4400
ALLPIS = 207'b001100011100000010100000110111010011000100101101011101010101101100001010100001111110001100010101001110111010110110010001110100111010110100111111101100111011101000101110111110000101101000000011010011110001000;
XPCT = 108'b001111110010110100000001101011110001100001111010101110010000001000011110111010100000101010011111000000100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4600

pattern = 23; // 4600
ALLPIS = 207'b111010111001110011011000001011111101111101011101010011110111010100001101111001010101010101011010101000111010011110111000100000101110001101010000011110101111110111000111000010010101111000100011001101111100011;
XPCT = 108'b111000010010111100010001100101111100011111111111011011001111111000010101000101011101111000000110100010001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4800

pattern = 24; // 4800
ALLPIS = 207'b100001101011001011100100010101101010100001100101010100100110001000001110010101000000111001111101011011111010001010101100001010100100010001100111100111100101111000110011111100011101110000110011000010111010110;
XPCT = 108'b111111100110111000011001100010111010111001011101111111101111010101001101111101001000110000000111010100010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5000

pattern = 25; // 5000
ALLPIS = 207'b110000110101100101110010001010110101010000110010101010010011000100000111001010100000011100111110101101111101000101010110000101010010001000110011110011110010111100011001111110001110111000011001100001011101011;
XPCT = 108'b110111110111011100001100110001011101110011111101111111101111100011101111100100110010111000100000110101010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5200

pattern = 26; // 5200
ALLPIS = 207'b000100101101000000110001010101001110110111010010101000010100000000001011001100111010011101001111011001011001100111011011011000011010010011010110010001001011011101011100100010010000010000101110010100101010010;
XPCT = 108'b000100010000001000010111001000101010101101110000101110011111011101101111111111011110111101000111100010000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5400

pattern = 27; // 5400
ALLPIS = 207'b100010010110100000011000101010100111011011101001010100001010000000000101100110011101001110100111101100101100110011101101101100001101001001101011001000100101101110101110010001001000001000010111001010010101001;
XPCT = 108'b111010000100000100001011100110010101000011111100001011101111100001001111010110101011111011000001001100001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5600

pattern = 28; // 5600
ALLPIS = 207'b001101111100100010000100000101000111110010111111010111011000100010001010011010100100110100000011111001110001011100000110101100110101110011111010001100100000110100000111010101110011001000101001000001001110011;
XPCT = 108'b001010101001100100010100100001001110111001110011111110010000111000000110000010001001101011111001010000110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5800

pattern = 29; // 5800
ALLPIS = 207'b100110111110010001000010000010100011111001011111101011101100010001000101001101010010011010000001111100111000101110000011010110011010111001111101000110010000011010000011101010111001100100010100100000100111001;
XPCT = 108'b111101011100110010001010010000100111011001111111011011111111010011011111000100010100110110000001101010000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6000

pattern = 30; // 6000
ALLPIS = 207'b110011011111001000100001000001010001111100101111110101110110001000100010100110101001001101000000111110011100010111000001101011001101011100111110100011001000001101000001110101011100110010001010010000010011100;
XPCT = 108'b110110100110011001000101001000010011011011111111011011101111100101111111010101011011110111011001011110100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6200

pattern = 31; // 6200
ALLPIS = 207'b111001101111100100010000100000101000111110010111111010111011000100010001010011010100100110100000011111001110001011100000110101100110101110011111010001100100000110100000111010101110011001000101001000001001110;
XPCT = 108'b110111011111001100100010100100001001100011111101111111001001111011011110011111011100110110000000001010000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6400

pattern = 32; // 6400
ALLPIS = 207'b001110011110000110111111000011100011111111010101000101000101001001100011010111101101110011110111100101111100001000101100001010011111101110100001101110101111101111100101000001010101110101011011111100101111001;
XPCT = 108'b000000000010111010101101111100101111011111111011011010000000110010011110001001111101100100011111111111110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6600

pattern = 33; // 6600
ALLPIS = 207'b111101111001100111010000110011011011000000100000010100010100011011111011100010010110101111001010011100100011001010100111001000111000010101001001110101000100010100011100010001000000101000001101000011100100111;
XPCT = 108'b110010000000010100000110100011100100100011111101111111101111100011101111011101101011111011011001110010000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6800

pattern = 34; // 6800
ALLPIS = 207'b000110001111011100010100101110100100110000110111100010100010101011101100000100111110100001111110110000001010111110010011111101011110011100100011000100101001011101010000100101101111000101110101010010000001100;
XPCT = 108'b000100101111100010111010101010000001000001111001011010011111110110001111110111011110110110111111010111111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7000

pattern = 35; // 7000
ALLPIS = 207'b100011000111101110001010010111010010011000011011110001010001010101110110000010011111010000111111011000000101011111001001111110101111001110010001100010010100101110101000010010110111100010111010101001000000110;
XPCT = 108'b110010011011110001011101010101000000001011110110000001001111011111011111101100000011111000100111111010110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7200

pattern = 36; // 7200
ALLPIS = 207'b111111111101110001111010001000001010110011011000111101101101100011011000010110100010011011101000001001111110100111001000110101001000001001101001011111100101111000110001001000001110000100000110101000001111010;
XPCT = 108'b110001000111000010000011010100001111010011111111011011111001111100011110100110100101110111111001111011010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7400

pattern = 37; // 7400
ALLPIS = 207'b011111111110111000111101000100000101011001101100011110110110110001101100001011010001001101110100000100111111010011100100011010100100000100110100101111110010111100011000100100000111000010000011010100000111101;
XPCT = 108'b000100100011100001000001101000000111000111111001011010000000110000001110011000111110101111111111110010011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7600

pattern = 38; // 7600
ALLPIS = 207'b000001100001011010100001100001100001010011100011001010011110010001010101010010000101010101001101100111100011100001011110000111001101101100111011111001010110110001101001010011010110010100011010010110101100111;
XPCT = 108'b000010010011001010001101001010101100111101111000101110001111101100010111111111101110111101000000100110001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7800

pattern = 39; // 7800
ALLPIS = 207'b100000110000101101010000110000110000101001110001100101001111001000101010101001000010101010100110110011110001110000101111000011100110110110011101111100101011011000110100101001101011001010001101001011010110011;
XPCT = 108'b110101001101100101000110100111010110100001111111111111101111101001011111011111110100111010000000001111011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8000

pattern = 40; // 8000
ALLPIS = 207'b010000011000010110101000011000011000010100111000110010100111100100010101010100100001010101010011011001111000111000010111100001110011011011001110111110010101101100011010010100110101100101000110100101101011001;
XPCT = 108'b001010101010110010100011010001101011101111011001111110001111001011110101010100001011110110000001011011011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8200

pattern = 41; // 8200
ALLPIS = 207'b100110010010001101101011001111101111110101001001011100010110111011101001111101111101011001011110001001000000010100100111111010100110000011000110110001100101011001101000001011001111000111111000101110011010101;
XPCT = 108'b110001010111100011111100010110011010000111111100001011111111101001101111111111110111110110000000110100001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8400

pattern = 42; // 8400
ALLPIS = 207'b111101010111000000001010100100010100000101110001101011001110010100010111101001010011011111011000100001011100000010111111110111001100101111000010110110011101000011010001000100110010010110100111101011100010011;
XPCT = 108'b110000101001001011010011110111100010111011111111111111111001100111001110001111111101110101100111110011011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8600

pattern = 43; // 8600
ALLPIS = 207'b011110101011100000000101010010001010000010111000110101100111001010001011110100101001101111101100010000101110000001011111111011100110010111100001011011001110100001101000100010011001001011010011110101110001001;
XPCT = 108'b000100010100100101101001111001110001001111111011011010011111001010111111110111001100111011011000111100011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8800

pattern = 44; // 8800
ALLPIS = 207'b000001001011110110111101101010100110111110001001011111110110101100100110101101111001000100000001101101101011001000000011110111101100100101010001000011001000111111010001010000011001010000110010000110010111101;
XPCT = 108'b000010000100101000011001000010010111111111111011111110001111110000101111100111111111110100111001001010110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9000

pattern = 45; // 9000
ALLPIS = 207'b000000100101111011011110110101010011011111000100101111111011010110010011010110111100100010000000110110110101100100000001111011110110010010101000100001100100011111101000101000001100101000011001000011001011110;
XPCT = 108'b000101000110010100001100100011001011100011111010101110011111011011000101111101100100111010111110110110101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9200

pattern = 46; // 9200
ALLPIS = 207'b001110001100111011010000011001001010010000110111010010111000100010101010111100110011100010110111111110100110111010101100110111100100100111110101111110011101100000010001010101010011100001010111011101001010110;
XPCT = 108'b000010100001110000101011101101001010011101101001011010000000111101100100001010001011101110011000111010111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9400

pattern = 47; // 9400
ALLPIS = 207'b101001011000011011010111001111000110110111001110101100011001011000110110001001110100000010101100011010101111010101111010010001101101111101011011010001100001011111101101101011111100000101110000010010001010010;
XPCT = 108'b110101011110000010111000001010001010111001111100100101010000101111011110011000011011101111000110000100000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9600

pattern = 48; // 9600
ALLPIS = 207'b011010010110000110110101110011110001101101110011101011000110010110001101100010011101000000101011000110101011110101011110100100011011011111010110110100011000010111111011011010111111000001011100000100100010100;
XPCT = 108'b001011011111100000101110000000100010011111111011011010011111101101011111001100000001111111000001101101010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9800

pattern = 49; // 9800
ALLPIS = 207'b001101001011000011011010111001111000110110111001110101100011001011000110110001001110100000010101100011010101111010101111010010001101101111101011011010001100001011111101101101011111100000101110000010010001010;
XPCT = 108'b000101100111110000010111000010010001111011111010101110011111110111101111101101100100111110000110001010111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10000

pattern = 50; // 10000
ALLPIS = 207'b111101001100110110001001101101111101110010111011011000011101111011010010111011111110011011110010111101001001010110000111111110111100110101011011011000001100101101011010011010000010001101010000011100001011011;
XPCT = 108'b111011010001000110101000001100001011100111111101111111110000101010100100110000100011100100100110111000001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10200

pattern = 51; // 10200
ALLPIS = 207'b100110000010001000000010111001001101011100010001010001100000110011100110010010100100101100110000111000010000011001011011110000111111010100100111101111111011010011000001000111011111101100100010000101111010011;
XPCT = 108'b110000110111110110010001000001111010011101111111011011110000111000011110101010011101100001000111100001111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10400

pattern = 52; // 10400
ALLPIS = 207'b010011000001000100000001011100100110101110001000101000110000011001110011001001010010010110011000011100001000001100101101111000011111101010010011110111111101101001100000100011101111110110010001000010111101001;
XPCT = 108'b000100011111111011001000100010111101000011111001011010011111011001001111100100111000111001011111010001100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10600

pattern = 53; // 10600
ALLPIS = 207'b100111111110100100111111101101110000101000010001010001011101000101011010110011000100111000111011101011111000001110111010110110010000011011101000010101010001011011010101010000100010001110010011011101110001101;
XPCT = 108'b110010001001000111001001101101110001010111111111011011101111100110101111101111110111111111100000110100000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10800

pattern = 54; // 10800
ALLPIS = 207'b100111100001101111110000111000111111110101010001010001010010011000110101111011011100111101111001011111000010001011000010100111111011101000011011101011111011111001010000010101011101010110111111001011110011010;
XPCT = 108'b110010100110101011011111100111110011001001111111010001111111100110111111010100011011110011100111100000100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11000

pattern = 55; // 11000
ALLPIS = 207'b110011110000110111111000011100011111111010101000101000101001001100011010111101101110011110111100101111100001000101100001010011111101110100001101110101111101111100101000001010101110101011011111100101111001101;
XPCT = 108'b110001011111010101101111110001111001000111011101011011100000111011111110010001111000100001111110110110111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11200

pattern = 56; // 11200
ALLPIS = 207'b111001111000011011111100001110001111111101010100010100010100100110001101011110110111001111011110010111110000100010110000101001111110111010000110111010111110111110010100000101010111010101101111110010111100110;
XPCT = 108'b110000100011101010110111111010111100101011011101111111100110000111001111011010011000100000111111100011111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11400

pattern = 57; // 11400
ALLPIS = 207'b011100111100001101111110000111000111111110101010001010001010010011000110101111011011100111101111001011111000010001011000010100111111011101000011011101011111011111001010000010101011101010110111111001011110011;
XPCT = 108'b001000011101110101011011111101011110100011111001111110010000001101001110111001001111101010000111111011011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11600

pattern = 58; // 11600
ALLPIS = 207'b101011111111011011101110000100010000001001101011010100001111110110010110000111011000100100100100011000001000100010000011110011100010110010001101111111101011010010001001101101111111011000001010100010110001111;
XPCT = 108'b110101101111101100000101010010110001011011111100001011001111111001111111000110001111110110100110010111100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11800

pattern = 59; // 11800
ALLPIS = 207'b110101111111101101110111000010001000000100110101101010000111111011001011000011101100010010010010001100000100010001000001111001110001011001000110111111110101101001000100110110111111101100000101010001011000111;
XPCT = 108'b110110111111110110000010101001011000101011111101111111000110000111001111101011001111100000111110100101001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12000

pattern = 60; // 12000
ALLPIS = 207'b110001000000101101010101100101010100001011110001100001001100001011110011100110101110101101101101011110001010101010100011001111011010011110101110100000010001100110101011110110100000101110001000001010011101100;
XPCT = 108'b111110111000010111000100000110011101110011111111111111101111001001101111100111010010111101100000111111000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12200

pattern = 61; // 12200
ALLPIS = 207'b010011011111001101000100110110111010001100010011100100101001110011101111110100001111110010010010110111001101110111010010010100001111111101011010101111100011100001011100010110101111001111001110100111111111001;
XPCT = 108'b000010111111100111100111010011111111000111111001011010011111010010001111100111110001110011011110000101100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12400

pattern = 62; // 12400
ALLPIS = 207'b010001001000011110100110001111100110100111110001010011001101100111110000111110101111101110110110100001110111001100110101011100110010100110010000010100001101010001010011110011010100011111110110111000100111001;
XPCT = 108'b001110010010001111111011011100100111111011111011111110011001010101111100110111000001111100100001111001001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12600

pattern = 63; // 12600
ALLPIS = 207'b100011011011010100111101000011100011011010010011111101101001000101101110011000001111010011111111001000110011000100011001011101111011100001000101110101101101111010100000010100010101010111110001111110100010011;
XPCT = 108'b110010100010101011111000111110100010001111110111011011011111011010011011000101011110110110000111111001011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12800

pattern = 64; // 12800
ALLPIS = 207'b010001101101101010011110100001110001101101001001111110110100100010110111001100000111101001111111100100011001100010001100101110111101110000100010111010110110111101010000001010001010101011111000111111010001001;
XPCT = 108'b000001010101010101111100011111010001100111111001111110011111010111111111101100101010111011011001110001000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13000

pattern = 65; // 13000
ALLPIS = 207'b110000110010011011101000010101001010001111110011111010110101011001110011011000010110110100000110111010100001000100110001011001001111000010100111001000101100000011001000011010001110100011011101101111010110010;
XPCT = 108'b110011010111010001101110110111010110100111111101111111000000111110100100011000110011101110111000011001101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13200

pattern = 66; // 13200
ALLPIS = 207'b010011100110010110011010001110110101001110010010101001010101011010101111101011010011111110100111000101011000000000011011011111000101010011011110011011111101010011101101100000111000001001100100010101011010110;
XPCT = 108'b000100001100000100110010001001011010011111111011011010001001101011001110010100101001111001100000000010000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13400

pattern = 67; // 13400
ALLPIS = 207'b000010001100010000100011000011001010101110100010000000100101011011000001110010110001011011110111111010100100100010001110011100000000011011100010110010010101111011111111011101100011011100111000101000011100100;
XPCT = 108'b001011101001101110011100010100011100010001111000001010001111101011101111100111100011110000000001100011011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13600

pattern = 68; // 13600
ALLPIS = 207'b011011011100011111100110110100100010100010000011110100000110100000100110011011110100110010011001100110100001101010100000010100100010110100110101010011001110001100110110011010100111101111000100101000110110110;
XPCT = 108'b001011011011110111100010010100110110000011111001011010000000010001001110011001100111100001000110111111000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13800

pattern = 69; // 13800
ALLPIS = 207'b110101011011010101100101110000111100011001001110100000101000111001011001110111101010010000100101011000111000111110010110001000110111111101101101101010000111001010101011101000010100001001110111010110101111110;
XPCT = 108'b111101000010000100111011101010101111111111010101111111001001111100000110000101111101111010011000101011101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14000

pattern = 70; // 14000
ALLPIS = 207'b011010101101101010110010111000011110001100100111010000010100011100101100111011110101001000010010101100011100011111001011000100011011111110110110110101000011100101010101110100001010000100111011101011010111111;
XPCT = 108'b000110100101000010011101110111010111010011111001011010011111111011001111001110001010110111011000011010010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14200

pattern = 71; // 14200
ALLPIS = 207'b101101010110110101011001011100001111000110010011101000001010001110010110011101111010100100001001010110001110001111100101100010001101111111011011011010100001110010101010111010000101000010011101110101101011111;
XPCT = 108'b111111010010100001001110111001101011100111111100101111000000010010000110111010000010101111100110011000010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14400

pattern = 72; // 14400
ALLPIS = 207'b010110101011011010101100101110000111100011001001110100000101000111001011001110111101010010000100101011000111000111110010110001000110111111101101101101010000111001010101011101000010100001001110111010110101111;
XPCT = 108'b000011100001010000100111011110110101010011111001011010011111100000011111100110010011111110011001101011010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14600

pattern = 73; // 14600
ALLPIS = 207'b001011010101101101010110010111000011110001100100111010000010100011100101100111011110101001000010010101100011100011111001011000100011011111110110110110101000011100101010101110100001010000100111011101011010111;
XPCT = 108'b001101111000101000010011101101011010000101111000001010001001001101101110001101100110111011000001011010101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14800

pattern = 74; // 14800
ALLPIS = 207'b101101100101101101001000010101100100010001001000101100011011100100100100001001111001001010110111000000100010100111111101111101101111011100010110101001010001001100001010010101101011001000001001100000101110001;
XPCT = 108'b111010101101100100000100110000101110100011111100101111111111011111101111111101001011111011111000100001100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15000

pattern = 75; // 15000
ALLPIS = 207'b101000010011000000011110000000100100100110111100101111100100100111101111100010100011011011000100110100000000000101111110010110011100100010100100001010111111100000100101100100010010110101000100011101011101001;
XPCT = 108'b110100100001011010100010001101011101111111111111111111101111000101111111100110101100110100111110110010111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15200

pattern = 76; // 15200
ALLPIS = 207'b101111111101101110111000010001000000100110101101010000111111011001011000011101100010010010010001100000100010001000001111001110001011001000110111111110101101001000100110110111111101100000101010001011000111110;
XPCT = 108'b111110111110110000010101000111000111001011111101011011000110001100111101010001111010101110011111011000110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15400

pattern = 77; // 15400
ALLPIS = 207'b010111111110110111011100001000100000010011010110101000011111101100101100001110110001001001001000110000010001000100000111100111000101100100011011111111010110100100010011011011111110110000010101000101100011111;
XPCT = 108'b001011011111011000001010100001100011011111111001011010000000101001110010000010100101100111000111001001100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15600

pattern = 78; // 15600
ALLPIS = 207'b110110100111000110110110011100110010001111101100110011010110101111000011101101110000111110001010100001011011110100100100100000111111101001100001111110001111000110010010010001000111100010001111011010111011100;
XPCT = 108'b111010000011110001000111101110111011000011111111011011101111000011001111011111001001111101111111000100100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15800

pattern = 79; // 15800
ALLPIS = 207'b010110011101101110110111110111111101011000101111111111000110001001100110101101011001100011010000010010011010010011011011010001100000100111110011000011011001101111101101101010101100110101011001011000101010110;
XPCT = 108'b000101011110011010101100101100101010010011111011011010001111010111111111101101100100110100100111010100111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16000

pattern = 80; // 16000
ALLPIS = 207'b011010101101101001100001001111101110001110110110001100001111111010110000001100110000001010111111111011000101000111011111110100101001011111110100010000110111111000110111111000010111111110101111001011100110100;
XPCT = 108'b001111000011111111010111100111100110011011011001011010011111100001100101110110010001111111111110110010001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16200

pattern = 81; // 16200
ALLPIS = 207'b101101010110110100110000100111110111000111011011000110000111111101011000000110011000000101011111111101100010100011101111111010010100101111111010001000011011111100011011111100001011111111010111100101110011010;
XPCT = 108'b111111100101111111101011110001110011110101111100101111010000000110001110101000100010100000011001010101111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16400

pattern = 82; // 16400
ALLPIS = 207'b011011100101010111110100101010011111111100110100000101101110100000101011011000101101111110111010111100000110111000111110111100110101000100111110111000010011110010101001011100001010111011110101000111001110101;
XPCT = 108'b000011100101011101111010100011001110010111101011011010001111011111001111100110000100111011011000101010001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16600

pattern = 83; // 16600
ALLPIS = 207'b110110111001010101111101001010100111111111001101000001011011101000001010110110001011011111101110101111000001101110001111101111001101010001001111101110000100111100101010010111000010101110111101010001110011101;
XPCT = 108'b111010110001010111011110101001110011000011011111011011101111100001011111010110001001110010111110101011110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16800

pattern = 84; // 16800
ALLPIS = 207'b011011000011101111000010111011111111110111100011000010110110100101100011001101111001111010110010000100001110000011000111001101011001110111011000111100111000000010111110001011011100000110111111011101101000001;
XPCT = 108'b001001010110000011011111101101101000001111111001011010011111001001001101001101100101111111111110101001011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17000

pattern = 85; // 17000
ALLPIS = 207'b100000101111111010001101100100011011100100101000000111110110001100110110111101011101000001001100000000110000101000101010100111010011101000101111100010000010001101111011100111100001000111000001011011000011000;
XPCT = 108'b111100111000100011100000101111000011110011111110100101011111110000101011000100011100110111011111001011111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17200

pattern = 86; // 17200
ALLPIS = 207'b010000010111111101000110110010001101110010010100000011111011000110011011011110101110100000100110000000011000010100010101010011101001110100010111110001000001000110111101110011110000100011100000101101100001100;
XPCT = 108'b000110011000010001110000010101100001111111111011111110001111100100101111001111011000111110111110001111110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17400

pattern = 87; // 17400
ALLPIS = 207'b101111101100110100001011001001110101001100010000010101000101000000100010000001111010101010010110000011101010011000101000110101111010100111100111111110000001011011011001101111110100101110101001100100010100111;
XPCT = 108'b110101111010010111010100110000010100011111111110001011100000011011111110101011110100100010000000101110110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17600

pattern = 88; // 17600
ALLPIS = 207'b101011111011001101000010110010011101010011000100000101010001010000001000100000011110101010100101100000111010100110001010001101011110101001111001111111100000010110110110011011111101001011101010011001000101001;
XPCT = 108'b111011011110100101110101001101000101001001111111011011111111000010001111000100101001111101011001101110110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17800

pattern = 89; // 17800
ALLPIS = 207'b111010111110110011010000101100100111010100110001000001010100010100000010001000000111101010101001011000001110101001100010100011010111101010011110011111111000000101101101100110111111010010111010100110010001010;
XPCT = 108'b110100111111101001011101010010010001011111111111011011100000000011111010000010001100101100100110110101000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18000

pattern = 90; // 18000
ALLPIS = 207'b010000010001010100000100101111110111110101000001000110000111010100000110011111100010001001000001101110110000111101111000010000010100100110001100110011100010001110010010010001010000101101000011100110111111101;
XPCT = 108'b001010000000010110100001110010111111101111111001111110011111100101010101011110001011110010011110011110011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18200

pattern = 91; // 18200
ALLPIS = 207'b100101000110100111101110101110011111100101111001000101101110110100000100010100010000111000110101110101101111110111110101001001110101000000000101100101101111001011101101101010100111010010111111000110101000110;
XPCT = 108'b110101011011101001011111100010101000110111100110101111100000110010001110001000100100101110100111111010011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18400

pattern = 92; // 18400
ALLPIS = 207'b101111110110101111001101110111010101110110110010100010001101000010000010101000110100110000000111111100000000001001011001110010100010111001100000100111010100110100101001001011101110010110100000101011010001101;
XPCT = 108'b110001011111001011010000010111010001010011111100001011000000001111111110000011010111100101111111011100100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18600

pattern = 93; // 18600
ALLPIS = 207'b111101011010101101000101000001000111010010000000011011110101111111100011000111111101110010001011011110011011110110110010111100010111000111111001110111111010001011011000000011111100000111100111010000001111111;
XPCT = 108'b110000011110000011110011101000001111101011110111111111000000001011011110010000011101101000000110111100010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18800

pattern = 94; // 18800
ALLPIS = 207'b101001110001101101100111001100100011111011001100110101101011110000111011011100001111100010101000010110111101001001001000001111111010011000011111100011110001100100100100010001111000100011110110101110111000011;
XPCT = 108'b110010001100010001111011010110111000101101111111110101011111100000001111011111101010111111011000110110001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19000

pattern = 95; // 19000
ALLPIS = 207'b110100111000110110110011100110010001111101100110011010110101111000011101101110000111110001010100001011011110100100100100000111111101001100001111110001111000110010010010001000111100010001111011010111011100001;
XPCT = 108'b111001001110001000111101101011011100101111111101111111011111011101011011010111000111111101100001011000001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19200

pattern = 96; // 19200
ALLPIS = 207'b011010011100011011011001110011001000111110110011001101011010111100001110110111000011111000101010000101101111010010010010000011111110100110000111111000111100011001001001000100011110001000111101101011101110000;
XPCT = 108'b000000100111000100011110110111101110011011111011011010011111001101010101001101101101111011100000110001100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19400

pattern = 97; // 19400
ALLPIS = 207'b001111101001101011100000000000110011100111000101110100011010111000000111111011100110000111011011011110010101100000100001001100101110011110011001101001101111111110101101011100100100010010011010010111010111101;
XPCT = 108'b000011101010001001001101001011010111010101111000001010001111100001101111000101000011111110011001110011110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19600

pattern = 98; // 19600
ALLPIS = 207'b010011000000100110011000000001011000010000111111000001101001100110001001110010010011101000011011010101011011111001101011000110111001000101001100100000101011111100011100110010100101110010001000011100001101001;
XPCT = 108'b000110011010111001000100001100001101000111111011011010010000011101111110100010001101100101011110000011110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19800

pattern = 99; // 19800
ALLPIS = 207'b101111111110010111010000011000111101001000111000000001001100010100000000010011000011101101011000011111011100110101010010110000010001111001000011011001110010010101000000100010101101100010000111010011100011000;
XPCT = 108'b110100011110110001000011101011100011000001111111011011110000110011011010010010001100101110111110001000110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20000

pattern = 100; // 20000
ALLPIS = 207'b010111111111001011101000001100011110100100011100000000100110001010000000001001100001110110101100001111101110011010101001011000001000111100100001101100111001001010100000010001010110110001000011101001110001100;
XPCT = 108'b000010000011011000100001110101110001001011111001011010001111101011011111111110101110110010111001101110110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20200

pattern = 101; // 20200
ALLPIS = 207'b100010100010100111001101000001001001100000000100101110010011010101010100000111011001001010000011010000100010100011100100100001111000010110110001010000111111001000101111110000111100101101011111000001110010010;
XPCT = 108'b111110001110010110101111100001110010011011111100001011111001110110011110100101011010110010100000011100011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20400

pattern = 102; // 20400
ALLPIS = 207'b010111000001000010010011010000100001111111000100111111111110001101010010111010010000010101111011101010011101001000011000000100110000011011110101111101100000001100100110100000101011011001001101100111001011001;
XPCT = 108'b001100001101101100100110110011001011000111111011011010011111111110010111000100111100110010011111001101001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20600

pattern = 103; // 20600
ALLPIS = 207'b101010100101010110000010011010101110011011011111101001101000010101101110010001000111000110011001101100001100111001110010101010011111010010001011110010110100000000011111000110110011000000011110110000000101000;
XPCT = 108'b111000111001100000001111011000000101011001111110001011011111010101111111000100001101111111011110001110010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20800

pattern = 104; // 20800
ALLPIS = 207'b011101010100101010110000010011010101110011011011111101001101000010101101110010001000111000110011001101100001100111001110010101010011111010010001011110010110100000000011111000110110011000000011110110000000101;
XPCT = 108'b001111001011001100000001111010000000111111111011111110000000000010111110101010010000101001011111100010101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21000

pattern = 105; // 21000
ALLPIS = 207'b010001111001000010011000001000001101110111100110010110010011010001011001001110001000010010101111011010011011110010100101010011110101000001111011111100010100101101011011000101010011101000110101010101101111001;
XPCT = 108'b001000100001110100011010101001101111111111111001111110011111000110001011010111000110110010111110101000000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21200

pattern = 106; // 21200
ALLPIS = 207'b110111101111110110001100000101100001110101111000100011111100011000100011010000001000000111100001010001100110111000010000110000100110011100001110101101010101101011110111011011100001010000101110000100011000111;
XPCT = 108'b111011011000101000010111000000011000010111101111011011001111111001001111000100000001111110000000101100100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21400

pattern = 107; // 21400
ALLPIS = 207'b100010010010010110000011000001101011111010011011111100100101111110001111001111100100000110100011001010001100001110100101000000100111111001011010000010111010100100010000101010011100000110010001110110010001100;
XPCT = 108'b110101010110000011001000111010010001001101111101011011001111000000001111111110110110110111000001110010000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21600

pattern = 108; // 21600
ALLPIS = 207'b010111001101001110000000110000101001011001100011001011010011100111100100001000011111000110110011101100110110100011001000011100100111100000001111001001000001010111101001010110000011010011111110001010110011110;
XPCT = 108'b000010110001101001111111000110110011010011111011011010000110100000111111010000111001101111111111100111110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21800

pattern = 109; // 21800
ALLPIS = 207'b111101001101011100000000000110011100111000101110100011010111000000111111011100110000111011011011110010101100000100001001100101110011110011001101001101111111110101101011100100100010010011010010111010111101101;
XPCT = 108'b111100101001001001101001011110111101110011011111111111101111001100101111000111001100111101111000000100100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22000

pattern = 110; // 22000
ALLPIS = 207'b011011001011100101110000010110011110110101010111111011000111110010001100111101010011010111101100001001011110101000101111000110001110010100011000101000011011110011100011000101111010101111101100110110101010000;
XPCT = 108'b001000101101010111110110011010101010011111111011011010011111010100101111100111011110110111011000011110101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22200

pattern = 111; // 22200
ALLPIS = 207'b000111100011110100011010111100100100110001110001001101000000101010110011000100001001110011010110101101001101110010110101101111011001100110001010000110100111011001110100111100110111010011011110011101001100100;
XPCT = 108'b000111101011101001101111001101001100001111111011010000001111101100111111101110101001111101011000100010110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22400

pattern = 112; // 22400
ALLPIS = 207'b010100110110001101010101111110110010101010110110010101011111011100000100111101110110011010010101011100100110011110001100110000000101011001011100010111001111100000011101111000100110010100100100111000001101101;
XPCT = 108'b000111001011001010010010011100001101110011011011111110001111110111111111001100110000110101000001110110011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22600

pattern = 113; // 22600
ALLPIS = 207'b001010011011000110101010111111011001010101011011001010101111101110000010011110111011001101001010101110010011001111000110011000000010101100101110001011100111110000001110111100010011001010010010011100000110110;
XPCT = 108'b001111100001100101001001001100000110001111111000001010001111100111011011111110110010111010011000100011110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22800

pattern = 114; // 22800
ALLPIS = 207'b000010100110110001101010101111110110010101010110110010101011111011100000100111101110110011010010101011100100110011110001100110000000101011001011100010111001111100000011101111000100110010100100100111000001101;
XPCT = 108'b001101110010011001010010010011000001010111111001011010011111001111111111101101100110111100100000010001101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23000

pattern = 115; // 23000
ALLPIS = 207'b100011011001110111110111000011100011000100111011110110011011111111101011100100100010101101001010001001010101010001011010010001110100110101011000100100000011010110111111000100000010110001111111001100100100010;
XPCT = 108'b111000100001011000111111100100100100010101111100001011111111011010011111011111100100111110011000000000010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23200

pattern = 116; // 23200
ALLPIS = 207'b110010001101110001101000100100101101010010110110101100111010100111111010001010011011001100100001010001010111001011001101111010000001101001010011101010100001111001111000000101010111000010110011110011011101010;
XPCT = 108'b110000100011100001011001111011011101001011111101011011101111111011110101010111011111111110111000101011011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23400

pattern = 117; // 23400
ALLPIS = 207'b110001001101111001000000001011110110101100000000110000100011111100110011100101100101111010111011100101110011101100100000111111111000111100000100000010101010000101001011111001010110101110000110110100001111001;
XPCT = 108'b111111000011010111000011011000001111111111110101111111111111110010101111010111100010111000011000001000110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23600

pattern = 118; // 23600
ALLPIS = 207'b011110101001011101100001111100111110111101101110010011010111011110001111100010110110111010101000101001110000001100111011111111101111001010011000100111111001000110010011000111110000111001101111111101000111110;
XPCT = 108'b001000111000011100110111111101000111011111111011011010010110111101101011101001101101101001111111011011000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23800

pattern = 119; // 23800
ALLPIS = 207'b110111110101000101011001101101111010111010100101111110100000001000101110110101000011001100010101100000000010100110011010110100111100000111010110100001110001101000011010100001001110110000011111110110101010111;
XPCT = 108'b111100000111011000001111111010101010000111111101011011101111101001101111001111001100110000011111011010011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24000

pattern = 120; // 24000
ALLPIS = 207'b010100011011000011100010100101101000000101110000110000100101111100100001011000001001011111111100110100101000101010001100110101000101100100000110010101111111011101000000100101011110111011010110011100001110101;
XPCT = 108'b000100100111011101101011001100001110101111111001111110011111100010101011110100101110111000111110101001001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24200

pattern = 121; // 24200
ALLPIS = 207'b011111010110100000100011001101001101010000000001110001000000100011101001010011000011110001110011110000011000111001100011101101011001101000110110101111111000011101000110000000101101001111101011100001011101111;
XPCT = 108'b001000001110100111110101110001011101000011111011011010000000100010100110110001111101100011111110100111111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24400

pattern = 122; // 24400
ALLPIS = 207'b100111110111100000011010010000011100101100100011001011011011011011000110000011101000111110101111011101011000010111010001001101111000000001101100111011010010000000101100011101000011011000111010000001001011000;
XPCT = 108'b110011100001101100011101000001001011000011110110001011111111100001101111100110111000110111111001001011001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24600

pattern = 123; // 24600
ALLPIS = 207'b110111010000111001000000111110011101101011001011010000110111110001100011000110111101101100001100010111100111110110110011001001101101010001110110010001000100011010000111000110001010101001011001100010101001000;
XPCT = 108'b111000110101010100101100110010101001010011001101011011111111001110110101111101110110110110100001011111110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24800

pattern = 124; // 24800
ALLPIS = 207'b100001111011000100101001100110101101111000001111010010101101101001110110011010000110010001000001100101101100101010010111110011001010111011001110100010100100111001110110100101000111011100110010101001111010001;
XPCT = 108'b111100100011101110011001010101111010100011111101110101011111010111101101101110001011111001011110100010010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25000

pattern = 125; // 25000
ALLPIS = 207'b111101011010000010001100110100110101000000000111000100000010001110100101001100001111000111001111000001100011100110001110110101100110100011011010111111100001110100011000000010110100111110101110000101110111100;
XPCT = 108'b110000011010011111010111000001110111101111111101111111000000011101011010110001001111100001011110001110100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25200

pattern = 126; // 25200
ALLPIS = 207'b111101110110111001111101011010010110101011111100101110101110111111010100100101101011111011011001100101101100101100111001001100000010011101101010000101001111001101000001010000110101011110000101101000011100101;
XPCT = 108'b110010001010101111000010110100011100111011110101111111100000010101101110101010001011100001111111101010000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25400

pattern = 127; // 25400
ALLPIS = 207'b011010111110101111100010101011010011110100010101001111100110001100100011001001100010100100100110110000101000011010000010110001111101111101101101011100101010010111111000101000000101000001101000010111001001101;
XPCT = 108'b000101000010100000110100001011001001000111111011011010001111101001000101011100000100111111100001001011011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25600

pattern = 128; // 25600
ALLPIS = 207'b110111000011010100110100000110101000111000011001001100000011101010010100111111111001101100100101000110101010010111110110011000110110010111100110110000000100100101111011010110000101010110100010011011111100011;
XPCT = 108'b111010110010101011010001001111111100010011011101011011111001001110011110111111111001110100100000000011110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25800

pattern = 129; // 25800
ALLPIS = 207'b101010001011111011111110110010000100101000011000000111001000011111101010010011110101001000111001000110100001010010101101101011011101101010000110110100100011011101111001101000011000110110011011000011000001101;
XPCT = 108'b110101000100011011001101100011000001011011111110001011111111001111001111000110100100110100111111001100100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26000

pattern = 130; // 26000
ALLPIS = 207'b001110010010010110111011000011111011000111110110100010011100100001110001101010101001101011110111100000111000100001101010100101101110111010001111111101001000011100001101110111110011100110101111111111000101101;
XPCT = 108'b000110111001110011010111111111000101011111111000000000000000110100011110000001101010100110011111100001011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26200

pattern = 131; // 26200
ALLPIS = 207'b000101011110010010000111110100000110000010111010010001110001101011000000010001100100110110110011011111111100010001100001000100011110110110101010011011111111000111011101100001101000100100001010010111000011100;
XPCT = 108'b000100001100010010000101001011000011110101111010101110001111001100111111110100100110111101000001000110100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26400

pattern = 132; // 26400
ALLPIS = 207'b010001111101011110001100010100011011101000100000010101011010100001010111110010010111000110101110101000011101000100101011011110000100001110010000101010100010001101000100101011001100011001001101011101010100001;
XPCT = 108'b000101010110001100100110101101010100100111111011111110011111000011101111101100111110110011011001111111101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26600

pattern = 133; // 26600
ALLPIS = 207'b001111010101101111010001111000011110111110011101110110101010011000100010010111100000001100111000110001011100010111111000001100011110111000000010000101010111110001100101000001101011100111010111100110100111010;
XPCT = 108'b000000001101110011101011110010100111010101111001011010011111011001111101101100101111110110111001111100110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26800

pattern = 134; // 26800
ALLPIS = 207'b110001001000110110001011010011001001110101011010100110000111101110100100111001111111011010000101000001000101001011101011000100010000001100010000101100110110111111000101000101101011001011000001010111111110001;
XPCT = 108'b110000101101100101100000101011111110110111111101111111111001111000011110011100100000110011100001100101000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27000

pattern = 135; // 27000
ALLPIS = 207'b001000011101011011101010100001010110111100011000101101001110000100000111111110101011111011010010001010110000111011100011001001000000100111001101011010101010110000111000100101000011010111110110010110111011110;
XPCT = 108'b000100100001101011111011001010111011100111111010101110011111011100101111011111111100110100111001011110001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27200

pattern = 136; // 27200
ALLPIS = 207'b011011101000001110010101010000101000010110011000111000001100110100110111010011001111110001111010001110100100010001011100101000101001110101001100111100111101001111110111011000010110011011111000111001100111101;
XPCT = 108'b001011000011001101111100011101100111011011111001011010000110100010001111000010001000100110011110110010100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27400

pattern = 137; // 27400
ALLPIS = 207'b111101101010001010010110101010111001100111100101000100000000010001101110110001000101101111010000001010010001101010010011100010000110110011011011001001100110100010111110100110001010000011010001001110111100101;
XPCT = 108'b111100110101000001101000100110111100100111111101111111100000000010001110001000001111100000011111100100011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27600

pattern = 138; // 27600
ALLPIS = 207'b000110010110011001000110111110110111000001000100010000101101100000110010010011100010010001011000011000110010010111010000100011010101011011000010100100010000000001001010111000000110100101001000011111000010110;
XPCT = 108'b001111000011010010100100001111000010000101111000000000011001110101111110110100010010110110000000110111111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27800

pattern = 139; // 27800
ALLPIS = 207'b010000011110111011100111010001001010010011000000100100010000011010000001110100110100001101111011110000100010010001111010000000110001111110010000010101111110011101111101001111100011011010110010101000010000011;
XPCT = 108'b000001111001101101011001010100010000110011111001111110000110000001011111101011100111101000100110100101101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28000

pattern = 140; // 28000
ALLPIS = 207'b111011110110010101011011111110000011111100110100101001011110011110010010011101001000001100100010000111010101100010010110010001000010111000100111100011010010111000110010010110100000011010000011001001100011101;
XPCT = 108'b111010111000001101000001100101100011000010111111011011100000100010000010100010001100101110011111101000101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28200

pattern = 141; // 28200
ALLPIS = 207'b011000001100001001111010111110110101111001101001000001010100001111010111010110100011100001110110100111101101010000110111000101100100110001100100111100110001110000000001000011110110111001011001101010101111000;
XPCT = 108'b000000011011011100101100110110101111111011111011111110001111101000001111001101001101111000000000111001110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28400

pattern = 142; // 28400
ALLPIS = 207'b110101111010001100111110001101101011001110000000011011101111111100100101011010100010111110001000111101110111000101010110101100111100111110010010000110100110101111001100100001110011100100000010110111101010111;
XPCT = 108'b110100001001110010000001011011101010101111111111111111101001111111011100010101100110110000000001110001010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28600

pattern = 143; // 28600
ALLPIS = 207'b110101100001011110111011100100101111001000110000001100111001000000010011110100000001000000111110010111001001010001101010111011111001011010101010111001111110000100000110100010101001110010010101011011100000101;
XPCT = 108'b111100011100111001001010101111100000100011111101111111001111101011010111011110001000111100011110010101101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28800

pattern = 144; // 28800
ALLPIS = 207'b001001111101011110010101001000100001010001100101010101101100011001100110100100101101111010101101110000110010010110001010001100011111110101011111001011000110101111011101101001001111100001100011111101010001011;
XPCT = 108'b000101000111110000110001111101010001110101010010101110011111110110111111000111101010110000111000000010000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29000

pattern = 145; // 29000
ALLPIS = 207'b001000001110011001001011010110111001101101001100111011101011011001011010110011001001110110110001110001100100100011111011101000101001000100100101001010100110011101001001111010011001011010110111110001010101010;
XPCT = 108'b000111010100101101011011111001010101111011111010101110010000110100011110100000100000101001011000101100110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29200

pattern = 146; // 29200
ALLPIS = 207'b100101010110110010011101101110010101110101011110110101011000011010011001110010000011110010010000001000000001100101011111011110100000011010000001000001011001001101110010100010001011000101001111011011111010001;
XPCT = 108'b111100010101100010100111101111111010100010111111111111011001000010011110111101010100111111100000001111001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29400

pattern = 147; // 29400
ALLPIS = 207'b111010110000100110101001010110100100111001111000010101100100111110010001111011001100100001100111101110001001101000001010001010111110001001001001000001001001110001010011000011001011011010000001010100010000110;
XPCT = 108'b111000010101101101000000101000010000010111111111011011010000011001001110100011011101101000011001110001101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29600

      $display("// %t : Simulation of %0d patterns completed with %0d errors\n", $time, pattern+1, nofails);
      if (verbose >=2) $finish(2);
      /* else */ $finish(0);
   end
endmodule
