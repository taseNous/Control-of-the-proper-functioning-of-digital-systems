// Verilog pattern output written by  TetraMAX (TM)  B-2008.09-SP2-i081128_181834 
// Date: Wed Jul  6 12:11:08 2011
// Module tested: c7552

//     Uncollapsed Stuck Fault Summary Report
// -----------------------------------------------
// fault class                     code   #faults
// ------------------------------  ----  ---------
// Detected                         DT       6827
// Possibly detected                PT          0
// Undetectable                     UD          0
// ATPG untestable                  AU          0
// Not detected                     ND         61
// -----------------------------------------------
// total faults                              6888
// test coverage                            99.11%
// -----------------------------------------------
// 
//            Pattern Summary Report
// -----------------------------------------------
// #internal patterns                         241
//     #basic_scan patterns                   241
// -----------------------------------------------
// 
// There are no rule fails
// There are no clocks
// There are no constraint ports
// There are no equivalent pins
// There are no net connections

`timescale 1 ns / 1 ns

//
// --- NOTE: Remove the comment to define 'tmax_iddq' to activate processing of IDDQ events
//     Or use '+define+tmax_iddq' on the verilog compile line
//
//`define tmax_iddq

module AAA_tmax_testbench_1_16 ;
   parameter NAMELENGTH = 200; // max length of names reported in fails
   integer nofails, bit, pattern, lastpattern;
   integer error_banner; // flag for tracking displayed error banner
   integer loads;        // number of load_unloads for current pattern
   integer patm1;        // pattern - 1
   integer patp1;        // pattern + lastpattern
   integer prev_pat;     // previous pattern number
   integer report_interval; // report pattern progress every Nth pattern
   integer verbose;      // message verbosity level
   parameter NINPUTS = 207, NOUTPUTS = 108;
   wire [0:NOUTPUTS-1] PO; reg [0:NOUTPUTS-1] ALLPOS, XPCT, MASK;
   reg [0:NINPUTS-1] PI, ALLPIS;
   reg [0:8*(NAMELENGTH-1)] POnames [0:NOUTPUTS-1];
   event IDDQ;

   wire N1;
   wire N5;
   wire N9;
   wire N12;
   wire N15;
   wire N18;
   wire N23;
   wire N26;
   wire N29;
   wire N32;
   wire N35;
   wire N38;
   wire N41;
   wire N44;
   wire N47;
   wire N50;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N69;
   wire N70;
   wire N73;
   wire N74;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N82;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N94;
   wire N97;
   wire N100;
   wire N103;
   wire N106;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N118;
   wire N121;
   wire N124;
   wire N127;
   wire N130;
   wire N133;
   wire N134;
   wire N135;
   wire N138;
   wire N141;
   wire N144;
   wire N147;
   wire N150;
   wire N151;
   wire N152;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N178;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire N185;
   wire N186;
   wire N187;
   wire N188;
   wire N189;
   wire N190;
   wire N191;
   wire N192;
   wire N193;
   wire N194;
   wire N195;
   wire N196;
   wire N197;
   wire N198;
   wire N199;
   wire N200;
   wire N201;
   wire N202;
   wire N203;
   wire N204;
   wire N205;
   wire N206;
   wire N207;
   wire N208;
   wire N209;
   wire N210;
   wire N211;
   wire N212;
   wire N213;
   wire N214;
   wire N215;
   wire N216;
   wire N217;
   wire N218;
   wire N219;
   wire N220;
   wire N221;
   wire N222;
   wire N223;
   wire N224;
   wire N225;
   wire N226;
   wire N227;
   wire N228;
   wire N229;
   wire N230;
   wire N231;
   wire N232;
   wire N233;
   wire N234;
   wire N235;
   wire N236;
   wire N237;
   wire N238;
   wire N239;
   wire N240;
   wire N242;
   wire N245;
   wire N248;
   wire N251;
   wire N254;
   wire N257;
   wire N260;
   wire N263;
   wire N267;
   wire N271;
   wire N274;
   wire N277;
   wire N280;
   wire N283;
   wire N286;
   wire N289;
   wire N293;
   wire N296;
   wire N299;
   wire N303;
   wire N307;
   wire N310;
   wire N313;
   wire N316;
   wire N319;
   wire N322;
   wire N325;
   wire N328;
   wire N331;
   wire N334;
   wire N337;
   wire N340;
   wire N343;
   wire N346;
   wire N349;
   wire N352;
   wire N355;
   wire N358;
   wire N361;
   wire N364;
   wire N367;
   wire N382;
   wire N241_I;
   wire N387;
   wire N388;
   wire N478;
   wire N482;
   wire N484;
   wire N486;
   wire N489;
   wire N492;
   wire N501;
   wire N505;
   wire N507;
   wire N509;
   wire N511;
   wire N513;
   wire N515;
   wire N517;
   wire N519;
   wire N535;
   wire N537;
   wire N539;
   wire N541;
   wire N543;
   wire N545;
   wire N547;
   wire N549;
   wire N551;
   wire N553;
   wire N556;
   wire N559;
   wire N561;
   wire N563;
   wire N565;
   wire N567;
   wire N569;
   wire N571;
   wire N573;
   wire N582;
   wire N643;
   wire N707;
   wire N813;
   wire N881;
   wire N882;
   wire N883;
   wire N884;
   wire N885;
   wire N889;
   wire N945;
   wire N1110;
   wire N1111;
   wire N1112;
   wire N1113;
   wire N1114;
   wire N1489;
   wire N1490;
   wire N1781;
   wire N10025;
   wire N10101;
   wire N10102;
   wire N10103;
   wire N10104;
   wire N10109;
   wire N10110;
   wire N10111;
   wire N10112;
   wire N10350;
   wire N10351;
   wire N10352;
   wire N10353;
   wire N10574;
   wire N10575;
   wire N10576;
   wire N10628;
   wire N10632;
   wire N10641;
   wire N10704;
   wire N10706;
   wire N10711;
   wire N10712;
   wire N10713;
   wire N10714;
   wire N10715;
   wire N10716;
   wire N10717;
   wire N10718;
   wire N10729;
   wire N10759;
   wire N10760;
   wire N10761;
   wire N10762;
   wire N10763;
   wire N10827;
   wire N10837;
   wire N10838;
   wire N10839;
   wire N10840;
   wire N10868;
   wire N10869;
   wire N10870;
   wire N10871;
   wire N10905;
   wire N10906;
   wire N10907;
   wire N10908;
   wire N11333;
   wire N11334;
   wire N11340;
   wire N11342;
   wire N241_O;

   // map PI[] vector to DUT inputs and bidis
   assign N1 = PI[0];
   assign N5 = PI[1];
   assign N9 = PI[2];
   assign N12 = PI[3];
   assign N15 = PI[4];
   assign N18 = PI[5];
   assign N23 = PI[6];
   assign N26 = PI[7];
   assign N29 = PI[8];
   assign N32 = PI[9];
   assign N35 = PI[10];
   assign N38 = PI[11];
   assign N41 = PI[12];
   assign N44 = PI[13];
   assign N47 = PI[14];
   assign N50 = PI[15];
   assign N53 = PI[16];
   assign N54 = PI[17];
   assign N55 = PI[18];
   assign N56 = PI[19];
   assign N57 = PI[20];
   assign N58 = PI[21];
   assign N59 = PI[22];
   assign N60 = PI[23];
   assign N61 = PI[24];
   assign N62 = PI[25];
   assign N63 = PI[26];
   assign N64 = PI[27];
   assign N65 = PI[28];
   assign N66 = PI[29];
   assign N69 = PI[30];
   assign N70 = PI[31];
   assign N73 = PI[32];
   assign N74 = PI[33];
   assign N75 = PI[34];
   assign N76 = PI[35];
   assign N77 = PI[36];
   assign N78 = PI[37];
   assign N79 = PI[38];
   assign N80 = PI[39];
   assign N81 = PI[40];
   assign N82 = PI[41];
   assign N83 = PI[42];
   assign N84 = PI[43];
   assign N85 = PI[44];
   assign N86 = PI[45];
   assign N87 = PI[46];
   assign N88 = PI[47];
   assign N89 = PI[48];
   assign N94 = PI[49];
   assign N97 = PI[50];
   assign N100 = PI[51];
   assign N103 = PI[52];
   assign N106 = PI[53];
   assign N109 = PI[54];
   assign N110 = PI[55];
   assign N111 = PI[56];
   assign N112 = PI[57];
   assign N113 = PI[58];
   assign N114 = PI[59];
   assign N115 = PI[60];
   assign N118 = PI[61];
   assign N121 = PI[62];
   assign N124 = PI[63];
   assign N127 = PI[64];
   assign N130 = PI[65];
   assign N133 = PI[66];
   assign N134 = PI[67];
   assign N135 = PI[68];
   assign N138 = PI[69];
   assign N141 = PI[70];
   assign N144 = PI[71];
   assign N147 = PI[72];
   assign N150 = PI[73];
   assign N151 = PI[74];
   assign N152 = PI[75];
   assign N153 = PI[76];
   assign N154 = PI[77];
   assign N155 = PI[78];
   assign N156 = PI[79];
   assign N157 = PI[80];
   assign N158 = PI[81];
   assign N159 = PI[82];
   assign N160 = PI[83];
   assign N161 = PI[84];
   assign N162 = PI[85];
   assign N163 = PI[86];
   assign N164 = PI[87];
   assign N165 = PI[88];
   assign N166 = PI[89];
   assign N167 = PI[90];
   assign N168 = PI[91];
   assign N169 = PI[92];
   assign N170 = PI[93];
   assign N171 = PI[94];
   assign N172 = PI[95];
   assign N173 = PI[96];
   assign N174 = PI[97];
   assign N175 = PI[98];
   assign N176 = PI[99];
   assign N177 = PI[100];
   assign N178 = PI[101];
   assign N179 = PI[102];
   assign N180 = PI[103];
   assign N181 = PI[104];
   assign N182 = PI[105];
   assign N183 = PI[106];
   assign N184 = PI[107];
   assign N185 = PI[108];
   assign N186 = PI[109];
   assign N187 = PI[110];
   assign N188 = PI[111];
   assign N189 = PI[112];
   assign N190 = PI[113];
   assign N191 = PI[114];
   assign N192 = PI[115];
   assign N193 = PI[116];
   assign N194 = PI[117];
   assign N195 = PI[118];
   assign N196 = PI[119];
   assign N197 = PI[120];
   assign N198 = PI[121];
   assign N199 = PI[122];
   assign N200 = PI[123];
   assign N201 = PI[124];
   assign N202 = PI[125];
   assign N203 = PI[126];
   assign N204 = PI[127];
   assign N205 = PI[128];
   assign N206 = PI[129];
   assign N207 = PI[130];
   assign N208 = PI[131];
   assign N209 = PI[132];
   assign N210 = PI[133];
   assign N211 = PI[134];
   assign N212 = PI[135];
   assign N213 = PI[136];
   assign N214 = PI[137];
   assign N215 = PI[138];
   assign N216 = PI[139];
   assign N217 = PI[140];
   assign N218 = PI[141];
   assign N219 = PI[142];
   assign N220 = PI[143];
   assign N221 = PI[144];
   assign N222 = PI[145];
   assign N223 = PI[146];
   assign N224 = PI[147];
   assign N225 = PI[148];
   assign N226 = PI[149];
   assign N227 = PI[150];
   assign N228 = PI[151];
   assign N229 = PI[152];
   assign N230 = PI[153];
   assign N231 = PI[154];
   assign N232 = PI[155];
   assign N233 = PI[156];
   assign N234 = PI[157];
   assign N235 = PI[158];
   assign N236 = PI[159];
   assign N237 = PI[160];
   assign N238 = PI[161];
   assign N239 = PI[162];
   assign N240 = PI[163];
   assign N242 = PI[164];
   assign N245 = PI[165];
   assign N248 = PI[166];
   assign N251 = PI[167];
   assign N254 = PI[168];
   assign N257 = PI[169];
   assign N260 = PI[170];
   assign N263 = PI[171];
   assign N267 = PI[172];
   assign N271 = PI[173];
   assign N274 = PI[174];
   assign N277 = PI[175];
   assign N280 = PI[176];
   assign N283 = PI[177];
   assign N286 = PI[178];
   assign N289 = PI[179];
   assign N293 = PI[180];
   assign N296 = PI[181];
   assign N299 = PI[182];
   assign N303 = PI[183];
   assign N307 = PI[184];
   assign N310 = PI[185];
   assign N313 = PI[186];
   assign N316 = PI[187];
   assign N319 = PI[188];
   assign N322 = PI[189];
   assign N325 = PI[190];
   assign N328 = PI[191];
   assign N331 = PI[192];
   assign N334 = PI[193];
   assign N337 = PI[194];
   assign N340 = PI[195];
   assign N343 = PI[196];
   assign N346 = PI[197];
   assign N349 = PI[198];
   assign N352 = PI[199];
   assign N355 = PI[200];
   assign N358 = PI[201];
   assign N361 = PI[202];
   assign N364 = PI[203];
   assign N367 = PI[204];
   assign N382 = PI[205];
   assign N241_I = PI[206];

   // map DUT outputs and bidis to PO[] vector
   assign
      PO[0] = N387 ,
      PO[1] = N388 ,
      PO[2] = N478 ,
      PO[3] = N482 ,
      PO[4] = N484 ,
      PO[5] = N486 ,
      PO[6] = N489 ,
      PO[7] = N492 ,
      PO[8] = N501 ,
      PO[9] = N505 ,
      PO[10] = N507 ,
      PO[11] = N509 ,
      PO[12] = N511 ,
      PO[13] = N513 ,
      PO[14] = N515 ,
      PO[15] = N517 ,
      PO[16] = N519 ,
      PO[17] = N535 ,
      PO[18] = N537 ,
      PO[19] = N539 ,
      PO[20] = N541 ,
      PO[21] = N543 ,
      PO[22] = N545 ,
      PO[23] = N547 ,
      PO[24] = N549 ,
      PO[25] = N551 ,
      PO[26] = N553 ,
      PO[27] = N556 ,
      PO[28] = N559 ,
      PO[29] = N561 ,
      PO[30] = N563 ,
      PO[31] = N565 ;
   assign
      PO[32] = N567 ,
      PO[33] = N569 ,
      PO[34] = N571 ,
      PO[35] = N573 ,
      PO[36] = N582 ,
      PO[37] = N643 ,
      PO[38] = N707 ,
      PO[39] = N813 ,
      PO[40] = N881 ,
      PO[41] = N882 ,
      PO[42] = N883 ,
      PO[43] = N884 ,
      PO[44] = N885 ,
      PO[45] = N889 ,
      PO[46] = N945 ,
      PO[47] = N1110 ,
      PO[48] = N1111 ,
      PO[49] = N1112 ,
      PO[50] = N1113 ,
      PO[51] = N1114 ,
      PO[52] = N1489 ,
      PO[53] = N1490 ,
      PO[54] = N1781 ,
      PO[55] = N10025 ,
      PO[56] = N10101 ,
      PO[57] = N10102 ,
      PO[58] = N10103 ,
      PO[59] = N10104 ,
      PO[60] = N10109 ,
      PO[61] = N10110 ,
      PO[62] = N10111 ,
      PO[63] = N10112 ;
   assign
      PO[64] = N10350 ,
      PO[65] = N10351 ,
      PO[66] = N10352 ,
      PO[67] = N10353 ,
      PO[68] = N10574 ,
      PO[69] = N10575 ,
      PO[70] = N10576 ,
      PO[71] = N10628 ,
      PO[72] = N10632 ,
      PO[73] = N10641 ,
      PO[74] = N10704 ,
      PO[75] = N10706 ,
      PO[76] = N10711 ,
      PO[77] = N10712 ,
      PO[78] = N10713 ,
      PO[79] = N10714 ,
      PO[80] = N10715 ,
      PO[81] = N10716 ,
      PO[82] = N10717 ,
      PO[83] = N10718 ,
      PO[84] = N10729 ,
      PO[85] = N10759 ,
      PO[86] = N10760 ,
      PO[87] = N10761 ,
      PO[88] = N10762 ,
      PO[89] = N10763 ,
      PO[90] = N10827 ,
      PO[91] = N10837 ,
      PO[92] = N10838 ,
      PO[93] = N10839 ,
      PO[94] = N10840 ,
      PO[95] = N10868 ;
   assign
      PO[96] = N10869 ,
      PO[97] = N10870 ,
      PO[98] = N10871 ,
      PO[99] = N10905 ,
      PO[100] = N10906 ,
      PO[101] = N10907 ,
      PO[102] = N10908 ,
      PO[103] = N11333 ,
      PO[104] = N11334 ,
      PO[105] = N11340 ,
      PO[106] = N11342 ,
      PO[107] = N241_O ;

   // instantiate the design into the testbench
   c7552 dut (
      .N1(N1),
      .N5(N5),
      .N9(N9),
      .N12(N12),
      .N15(N15),
      .N18(N18),
      .N23(N23),
      .N26(N26),
      .N29(N29),
      .N32(N32),
      .N35(N35),
      .N38(N38),
      .N41(N41),
      .N44(N44),
      .N47(N47),
      .N50(N50),
      .N53(N53),
      .N54(N54),
      .N55(N55),
      .N56(N56),
      .N57(N57),
      .N58(N58),
      .N59(N59),
      .N60(N60),
      .N61(N61),
      .N62(N62),
      .N63(N63),
      .N64(N64),
      .N65(N65),
      .N66(N66),
      .N69(N69),
      .N70(N70),
      .N73(N73),
      .N74(N74),
      .N75(N75),
      .N76(N76),
      .N77(N77),
      .N78(N78),
      .N79(N79),
      .N80(N80),
      .N81(N81),
      .N82(N82),
      .N83(N83),
      .N84(N84),
      .N85(N85),
      .N86(N86),
      .N87(N87),
      .N88(N88),
      .N89(N89),
      .N94(N94),
      .N97(N97),
      .N100(N100),
      .N103(N103),
      .N106(N106),
      .N109(N109),
      .N110(N110),
      .N111(N111),
      .N112(N112),
      .N113(N113),
      .N114(N114),
      .N115(N115),
      .N118(N118),
      .N121(N121),
      .N124(N124),
      .N127(N127),
      .N130(N130),
      .N133(N133),
      .N134(N134),
      .N135(N135),
      .N138(N138),
      .N141(N141),
      .N144(N144),
      .N147(N147),
      .N150(N150),
      .N151(N151),
      .N152(N152),
      .N153(N153),
      .N154(N154),
      .N155(N155),
      .N156(N156),
      .N157(N157),
      .N158(N158),
      .N159(N159),
      .N160(N160),
      .N161(N161),
      .N162(N162),
      .N163(N163),
      .N164(N164),
      .N165(N165),
      .N166(N166),
      .N167(N167),
      .N168(N168),
      .N169(N169),
      .N170(N170),
      .N171(N171),
      .N172(N172),
      .N173(N173),
      .N174(N174),
      .N175(N175),
      .N176(N176),
      .N177(N177),
      .N178(N178),
      .N179(N179),
      .N180(N180),
      .N181(N181),
      .N182(N182),
      .N183(N183),
      .N184(N184),
      .N185(N185),
      .N186(N186),
      .N187(N187),
      .N188(N188),
      .N189(N189),
      .N190(N190),
      .N191(N191),
      .N192(N192),
      .N193(N193),
      .N194(N194),
      .N195(N195),
      .N196(N196),
      .N197(N197),
      .N198(N198),
      .N199(N199),
      .N200(N200),
      .N201(N201),
      .N202(N202),
      .N203(N203),
      .N204(N204),
      .N205(N205),
      .N206(N206),
      .N207(N207),
      .N208(N208),
      .N209(N209),
      .N210(N210),
      .N211(N211),
      .N212(N212),
      .N213(N213),
      .N214(N214),
      .N215(N215),
      .N216(N216),
      .N217(N217),
      .N218(N218),
      .N219(N219),
      .N220(N220),
      .N221(N221),
      .N222(N222),
      .N223(N223),
      .N224(N224),
      .N225(N225),
      .N226(N226),
      .N227(N227),
      .N228(N228),
      .N229(N229),
      .N230(N230),
      .N231(N231),
      .N232(N232),
      .N233(N233),
      .N234(N234),
      .N235(N235),
      .N236(N236),
      .N237(N237),
      .N238(N238),
      .N239(N239),
      .N240(N240),
      .N242(N242),
      .N245(N245),
      .N248(N248),
      .N251(N251),
      .N254(N254),
      .N257(N257),
      .N260(N260),
      .N263(N263),
      .N267(N267),
      .N271(N271),
      .N274(N274),
      .N277(N277),
      .N280(N280),
      .N283(N283),
      .N286(N286),
      .N289(N289),
      .N293(N293),
      .N296(N296),
      .N299(N299),
      .N303(N303),
      .N307(N307),
      .N310(N310),
      .N313(N313),
      .N316(N316),
      .N319(N319),
      .N322(N322),
      .N325(N325),
      .N328(N328),
      .N331(N331),
      .N334(N334),
      .N337(N337),
      .N340(N340),
      .N343(N343),
      .N346(N346),
      .N349(N349),
      .N352(N352),
      .N355(N355),
      .N358(N358),
      .N361(N361),
      .N364(N364),
      .N367(N367),
      .N382(N382),
      .N241_I(N241_I),
      .N387(N387),
      .N388(N388),
      .N478(N478),
      .N482(N482),
      .N484(N484),
      .N486(N486),
      .N489(N489),
      .N492(N492),
      .N501(N501),
      .N505(N505),
      .N507(N507),
      .N509(N509),
      .N511(N511),
      .N513(N513),
      .N515(N515),
      .N517(N517),
      .N519(N519),
      .N535(N535),
      .N537(N537),
      .N539(N539),
      .N541(N541),
      .N543(N543),
      .N545(N545),
      .N547(N547),
      .N549(N549),
      .N551(N551),
      .N553(N553),
      .N556(N556),
      .N559(N559),
      .N561(N561),
      .N563(N563),
      .N565(N565),
      .N567(N567),
      .N569(N569),
      .N571(N571),
      .N573(N573),
      .N582(N582),
      .N643(N643),
      .N707(N707),
      .N813(N813),
      .N881(N881),
      .N882(N882),
      .N883(N883),
      .N884(N884),
      .N885(N885),
      .N889(N889),
      .N945(N945),
      .N1110(N1110),
      .N1111(N1111),
      .N1112(N1112),
      .N1113(N1113),
      .N1114(N1114),
      .N1489(N1489),
      .N1490(N1490),
      .N1781(N1781),
      .N10025(N10025),
      .N10101(N10101),
      .N10102(N10102),
      .N10103(N10103),
      .N10104(N10104),
      .N10109(N10109),
      .N10110(N10110),
      .N10111(N10111),
      .N10112(N10112),
      .N10350(N10350),
      .N10351(N10351),
      .N10352(N10352),
      .N10353(N10353),
      .N10574(N10574),
      .N10575(N10575),
      .N10576(N10576),
      .N10628(N10628),
      .N10632(N10632),
      .N10641(N10641),
      .N10704(N10704),
      .N10706(N10706),
      .N10711(N10711),
      .N10712(N10712),
      .N10713(N10713),
      .N10714(N10714),
      .N10715(N10715),
      .N10716(N10716),
      .N10717(N10717),
      .N10718(N10718),
      .N10729(N10729),
      .N10759(N10759),
      .N10760(N10760),
      .N10761(N10761),
      .N10762(N10762),
      .N10763(N10763),
      .N10827(N10827),
      .N10837(N10837),
      .N10838(N10838),
      .N10839(N10839),
      .N10840(N10840),
      .N10868(N10868),
      .N10869(N10869),
      .N10870(N10870),
      .N10871(N10871),
      .N10905(N10905),
      .N10906(N10906),
      .N10907(N10907),
      .N10908(N10908),
      .N11333(N11333),
      .N11334(N11334),
      .N11340(N11340),
      .N11342(N11342),
      .N241_O(N241_O)   );


   integer errshown;
   event measurePO;
   always @ measurePO begin
      if (((XPCT&MASK) !== (ALLPOS&MASK)) || (XPCT !== (~(~XPCT)))) begin
         errshown = 0;
         for (bit = 0; bit < NOUTPUTS; bit=bit + 1) begin
            if (MASK[bit]==1'b1) begin
               if (XPCT[bit] !== ALLPOS[bit]) begin
                  if (errshown==0) $display("\n// *** ERROR during capture pattern %0d, T=%t", pattern, $time);
                  $display("  %0d %0s (exp=%b, got=%b)", pattern, POnames[bit], XPCT[bit], ALLPOS[bit]);
                  nofails = nofails + 1; errshown = 1;
               end
            end
         end
      end
   end

   event forcePI_default_WFT;
   always @ forcePI_default_WFT begin
      PI = ALLPIS;
   end
   event measurePO_default_WFT;
   always @ measurePO_default_WFT begin
      #40;
      ALLPOS = PO;
      #0; #0 -> measurePO;
      `ifdef tmax_iddq
         #0; ->IDDQ;
      `endif
   end

   always @ IDDQ begin
   `ifdef tmax_iddq
      $ssi_iddq("strobe_try");
      $ssi_iddq("status drivers leaky AAA_tmax_testbench_1_16.leaky");
   `endif
   end

   event capture;
   always @ capture begin
      ->forcePI_default_WFT;
      #100; ->measurePO_default_WFT;
   end


   initial begin

      //
      // --- establish a default time format for %t
      //
      $timeformat(-9,2," ns",18);

      //
      // --- default verbosity to 2 but also allow user override by
      //     using '+define+tmax_msg=N' on verilog compile line.
      //
      `ifdef tmax_msg
         verbose = `tmax_msg ;
      `else
         verbose = 2 ;
      `endif

      //
      // --- default pattern reporting interval to 5 but also allow user
      //     override by using '+define+tmax_rpt=N' on verilog compile line.
      //
      `ifdef tmax_rpt
         report_interval = `tmax_rpt ;
      `else
         report_interval = 5 ;
      `endif

      //
      // --- support generating Extened VCD output by using
      //     '+define+tmax_vcde' on verilog compile line.
      //
      `ifdef tmax_vcde
         // extended VCD, see IEEE Verilog P1364.1-1999 Draft 2
         if (verbose >= 2) $display("// %t : opening Extended VCD output file", $time);
         $dumpports( dut, "sim_vcde.out");
      `endif

      //
      // --- IDDQ PLI initialization
      //     User may activite by using '+define+tmax_iddq' on verilog compile line.
      //     Or by defining `tmax_iddq in this file.
      //
      `ifdef tmax_iddq
         if (verbose >= 3) $display("// %t : Initializing IDDQ PLI", $time);
         $ssi_iddq("dut AAA_tmax_testbench_1_16.dut");
         $ssi_iddq("verb on");
         $ssi_iddq("cycle 0");
         //
         // --- User may select one of the following two methods for fault seeding:
         //     #1 faults seeded by PLI (default)
         //     #2 faults supplied in a file
         //     Comment out the unused lines as needed (precede with '//').
         //     Replace the 'FAULTLIST_FILE' string with the actual file pathname.
         //
         $ssi_iddq("seed SA AAA_tmax_testbench_1_16.dut");   // no file, faults seeded by PLI
         //
         // $ssi_iddq("scope AAA_tmax_testbench_1_16.dut");   // set scope for faults from a file
         // $ssi_iddq("read_tmax FAULTLIST_FILE"); // read faults from a file
         //
      `endif

      POnames[0] = "N387";
      POnames[1] = "N388";
      POnames[2] = "N478";
      POnames[3] = "N482";
      POnames[4] = "N484";
      POnames[5] = "N486";
      POnames[6] = "N489";
      POnames[7] = "N492";
      POnames[8] = "N501";
      POnames[9] = "N505";
      POnames[10] = "N507";
      POnames[11] = "N509";
      POnames[12] = "N511";
      POnames[13] = "N513";
      POnames[14] = "N515";
      POnames[15] = "N517";
      POnames[16] = "N519";
      POnames[17] = "N535";
      POnames[18] = "N537";
      POnames[19] = "N539";
      POnames[20] = "N541";
      POnames[21] = "N543";
      POnames[22] = "N545";
      POnames[23] = "N547";
      POnames[24] = "N549";
      POnames[25] = "N551";
      POnames[26] = "N553";
      POnames[27] = "N556";
      POnames[28] = "N559";
      POnames[29] = "N561";
      POnames[30] = "N563";
      POnames[31] = "N565";
      POnames[32] = "N567";
      POnames[33] = "N569";
      POnames[34] = "N571";
      POnames[35] = "N573";
      POnames[36] = "N582";
      POnames[37] = "N643";
      POnames[38] = "N707";
      POnames[39] = "N813";
      POnames[40] = "N881";
      POnames[41] = "N882";
      POnames[42] = "N883";
      POnames[43] = "N884";
      POnames[44] = "N885";
      POnames[45] = "N889";
      POnames[46] = "N945";
      POnames[47] = "N1110";
      POnames[48] = "N1111";
      POnames[49] = "N1112";
      POnames[50] = "N1113";
      POnames[51] = "N1114";
      POnames[52] = "N1489";
      POnames[53] = "N1490";
      POnames[54] = "N1781";
      POnames[55] = "N10025";
      POnames[56] = "N10101";
      POnames[57] = "N10102";
      POnames[58] = "N10103";
      POnames[59] = "N10104";
      POnames[60] = "N10109";
      POnames[61] = "N10110";
      POnames[62] = "N10111";
      POnames[63] = "N10112";
      POnames[64] = "N10350";
      POnames[65] = "N10351";
      POnames[66] = "N10352";
      POnames[67] = "N10353";
      POnames[68] = "N10574";
      POnames[69] = "N10575";
      POnames[70] = "N10576";
      POnames[71] = "N10628";
      POnames[72] = "N10632";
      POnames[73] = "N10641";
      POnames[74] = "N10704";
      POnames[75] = "N10706";
      POnames[76] = "N10711";
      POnames[77] = "N10712";
      POnames[78] = "N10713";
      POnames[79] = "N10714";
      POnames[80] = "N10715";
      POnames[81] = "N10716";
      POnames[82] = "N10717";
      POnames[83] = "N10718";
      POnames[84] = "N10729";
      POnames[85] = "N10759";
      POnames[86] = "N10760";
      POnames[87] = "N10761";
      POnames[88] = "N10762";
      POnames[89] = "N10763";
      POnames[90] = "N10827";
      POnames[91] = "N10837";
      POnames[92] = "N10838";
      POnames[93] = "N10839";
      POnames[94] = "N10840";
      POnames[95] = "N10868";
      POnames[96] = "N10869";
      POnames[97] = "N10870";
      POnames[98] = "N10871";
      POnames[99] = "N10905";
      POnames[100] = "N10906";
      POnames[101] = "N10907";
      POnames[102] = "N10908";
      POnames[103] = "N11333";
      POnames[104] = "N11334";
      POnames[105] = "N11340";
      POnames[106] = "N11342";
      POnames[107] = "N241_O";
      nofails = 0; pattern = -1; lastpattern = 0;
      prev_pat = -2; error_banner = -2;
      /*** No test setup procedure ***/


      /*** Non-scan test ***/

      if (verbose >= 1) $display("// %t : Begin patterns, first pattern = 0", $time);
pattern = 0; // 0
ALLPIS = 207'b001100001101110001011100101010111000010011000000100100110001110001110010100001110000101101100100011011011010111011111000100110001001111101110100101010011010100001001011011010000011011010001011010110010000010;
XPCT = 108'b001011010001101101000101101010010000110111111000100100001001110111011110100101000011111001100000110000111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 200

pattern = 1; // 200
ALLPIS = 207'b000110000110111000101110010101011100001001100000010010011000111000111001010000111000010110110010001101101101011101111100010011000100111110111010010101001101010000100101101101000001101101000101101011001000001;
XPCT = 108'b000101100000110110100010110111001000010011111001010000011111111110011111001101100110110010000001011101001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 400

pattern = 2; // 400
ALLPIS = 207'b001111001110101101001011100000010110010111110000101101111101101101101110001001101100100110111101011101101100010101000110101111101011100010101001100000111100001001011001101100100011101100101001100011110100010;
XPCT = 108'b000101101001110110010100110011110100010011111010001010010000001110101110101010000100100010011000001001101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 600

pattern = 3; // 600
ALLPIS = 207'b001011101010100111111001011010110011011000111000110010001111000111000101100101000110111110111010110101101100110001011011110001111100001100100000011010000100100101100111101100010010101100011111100111101010011;
XPCT = 108'b001101100001010110001111110011101010011111111001011010010000011010101110001000011000100111011000010110011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 800

pattern = 4; // 800
ALLPIS = 207'b001001111000100010100000000111100001111111011100111101110110010010010000010011010011110010111001000001101100100011010101011110110111111011100100100111011000110011111000101100001010001100000100100101100101011;
XPCT = 108'b000101100101000110000010010001100101100101111010101110010000101011101110111011010011100000011110000100010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1000

pattern = 5; // 1000
ALLPIS = 207'b100100111100010001010000000011110000111111101110011110111011001001001000001001101001111001011100100000110110010001101010101111011011111101110010010011101100011001111100010110000101000110000010010010110010101;
XPCT = 108'b110010110010100011000001001010110010100001111100101111101111111100001111010100101011110111000001010010111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1200

pattern = 6; // 1200
ALLPIS = 207'b011110010011111001110100101011000000001100110111101011101100010101010110100101000100010001001010001011000001110011001101110001100100000011001101100011101100101101110101010001000001111001001010011111001001000;
XPCT = 108'b000010000000111100100101001111001001010111111011011010011111010111001111100110011001111000111000101000010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1400

pattern = 7; // 1400
ALLPIS = 207'b001111001001111100111010010101100000000110011011110101110110001010101011010010100010001000100101000101100000111001100110111000110010000001100110110001110110010110111010101000100000111100100101001111100100100;
XPCT = 108'b001101001000011110010010100111100100000111111010001010001111110101100111011100100100110001111001001100010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1600

pattern = 8; // 1600
ALLPIS = 207'b101011101001001111000001100000001000010000001101011110001010110100100111001000100001101001110110111001101010100111001011111010010000111101000111110010100001101010010110001110010011000100011001110001100010000;
XPCT = 108'b111001110001100010001100111001100010001001111101011011111111001110001111001101011100111001111001011101010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1800

pattern = 9; // 1800
ALLPIS = 207'b010101110100100111100000110000000100001000000110101111000101011010010011100100010000110100111011011100110101010011100101111101001000011110100011111001010000110101001011000111001001100010001100111000110001000;
XPCT = 108'b001000110100110001000110011100110001110011111011111110011111100001101111001101110111111111100001100011000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2000

pattern = 10; // 2000
ALLPIS = 207'b101010111010010011110000011000000010000100000011010111100010101101001001110010001000011010011101101110011010101001110010111110100100001111010001111100101000011010100101100011100100110001000110011100011000100;
XPCT = 108'b110100011010011000100011001100011000010101111111011011111111011001001111000111001100111100100001101111111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2200

pattern = 11; // 2200
ALLPIS = 207'b011001010000111000100100100110111001010001000001001111000000100111010110011000110100100000101010101100010111101111000001111001011011111010011100010100001110101100011001101011110001000010101000011000011100000;
XPCT = 108'b000101011000100001010100001100011100111011111011111110010000011000101110101010111110100010111111100110100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2400

pattern = 12; // 2400
ALLPIS = 207'b000000100101101101001110111001100100111011100000000011010001100010011001101101101010111101110001001101010001001100011000011010100100000000111010100000011101110111000111101111111011111011011111011010011110010;
XPCT = 108'b001101111101111101101111101110011110111011110011111110011111110101101111001100010100111000100001110011010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2600

pattern = 13; // 2600
ALLPIS = 207'b100000010010110110100111011100110010011101110000000001101000110001001100110110110101011110111000100110101000100110001100001101010010000000011101010000001110111011100011110111111101111101101111101101001111001;
XPCT = 108'b111110111110111110110111110101001111111101111111111111111111010010011111101100011000110000100001101010110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2800

pattern = 14; // 2800
ALLPIS = 207'b111100000100101010001111000100100001011101111000100100000101101001010100111010101010000010111000001000001110101000111110100000100000111101111010000010011101111100111010100001111101100100111100100000110111110;
XPCT = 108'b111100001110110010011110010000110111101011111101111111010000000101001110110001011110100110011110000010001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3000

pattern = 15; // 3000
ALLPIS = 207'b011110000010010101000111100010010000101110111100010010000010110100101010011101010101000001011100000100000111010100011111010000010000011110111101000001001110111110011101010000111110110010011110010000011011111;
XPCT = 108'b000010001111011001001111001000011011011011011001011010000000101010101110000011001011101100011111010011110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3200

pattern = 16; // 3200
ALLPIS = 207'b000011001100111011111111011011110000000100011110101101110000101011100111101111011010001101001010011001011001010001110111001110000001110010101010001010111101111110000101110010011100000011000100011110011101101;
XPCT = 108'b000110010110000001100010001110011101011111111011011010001111011011111111100101100011111101100000000110111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3400

pattern = 17; // 3400
ALLPIS = 207'b001101101011101100100011000111000000010001001111110010001001100100000001010110011101101011000001010111110110010011000011000001001001000100100001101111000100011110001001100011001101011011101001011001011110100;
XPCT = 108'b000100010110101101110100101101011110110001111000101110001111100101111111101110011110111001111000100111101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3600

pattern = 18; // 3600
ALLPIS = 207'b100110110101110110010001100011100000001000100111111001000100110010000000101011001110110101100000101011111011001001100001100000100100100010010000110111100010001111000100110001100110101101110100101100101111010;
XPCT = 108'b110110001011010110111010010100101111000101111111011011011111101011011011011100101000110010111111110111011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3800

pattern = 19; // 3800
ALLPIS = 207'b110011011010111011001000110001110000000100010011111100100010011001000000010101100111011010110000010101111101100100110000110000010010010001001000011011110001000111100010011000110011010110111010010110010111101;
XPCT = 108'b111011001001101011011101001010010111001111111101011011100000000010111110010010100111101011111110001001101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4000

pattern = 20; // 4000
ALLPIS = 207'b011001101101011101100100011000111000000010001001111110010001001100100000001010110011101101011000001010111110110010011000011000001001001000100100001101111000100011110001001100011001101011011101001011001011110;
XPCT = 108'b000001100100110101101110100111001011111011101001111110001111010111111111110110011001110101100111001001101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4200

pattern = 21; // 4200
ALLPIS = 207'b101100110110101110110010001100011100000001000100111111001000100110010000000101011001110110101100000101011111011001001100001100000100100100010010000110111100010001111000100110001100110101101110100101100101111;
XPCT = 108'b110100110110011010110111010001100101100101111110101111000000000110011110110011001100100100100000100110110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4400

pattern = 22; // 4400
ALLPIS = 207'b111010010110100110000101101100110110010011100010111011010101100010111010100011011100010110110010011001110101010111011110100000001011101111111101101001000100101001110111001001000101000000111100000100100010101;
XPCT = 108'b111001000010100000011110000000100010010111111111011011011111101100011011100100100101111111100001110001011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4600

pattern = 23; // 4600
ALLPIS = 207'b010001000110100010011110011100100011011010110001111001011011000000101111110000011110100110111101010111100000010000010111110110001100001010001010011110111000110101110000111110100001111010010101010100000001000;
XPCT = 108'b000111111000111101001010101000000001100111111011111110010000101010001110010001101000101010111111101000111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4800

pattern = 24; // 4800
ALLPIS = 207'b000100101110100000010011100100101001111110011000011000011100010001100101011001111111111110111010110000101010110011110011011101001111111000110001100101000110111011110011000101010011100111000001111100010000110;
XPCT = 108'b001000100001110011100000111100010000111101111001111110000000010100111110100011101111100101111111010001011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5000

pattern = 25; // 5000
ALLPIS = 207'b100010010111010000001001110010010100111111001100001100001110001000110010101100111111111111011101011000010101011001111001101110100111111100011000110010100011011101111001100010101001110011100000111110001000011;
XPCT = 108'b110100011100111001110000011110001000010111111100000001101111000011001111101111111110111011000110011001011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5200

pattern = 26; // 5200
ALLPIS = 207'b111101000110011001011000010011110010001100100110100010110110110101101011110111101111010010001010110111010000010111000100010001011010000011111000110011001011001111110111101011010111100011111011001001010100011;
XPCT = 108'b111101010011110001111101100101010100111011111101111111010000011110011100101010000110101110100111001000000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5400

pattern = 27; // 5400
ALLPIS = 207'b011110100011001100101100001001111001000110010011010001011011011010110101111011110111101001000101011011101000001011100010001000101101000001111100011001100101100111111011110101101011110001111101100100101010001;
XPCT = 108'b001110101101111000111110110000101010010111111011011010001111010010111111100101101000111100111001001100001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5600

pattern = 28; // 5600
ALLPIS = 207'b000011011100010111001010101110000100110000001001001100011100011100101000011100001011011001000110110110101110111110001001100010011111011101001010100110101000010010110110100000110110100010110101100100000101010;
XPCT = 108'b001100001011010001011010110000000101001111101001011010011001011010101110010101010010111111100000101000011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5800

pattern = 29; // 5800
ALLPIS = 207'b100001101110001011100101010111000010011000000100100110001110001110010100001110000101101100100011011011010111011111000100110001001111101110100101010011010100001001011011010000011011010001011010110010000010101;
XPCT = 108'b111010000101101000101101011010000010111001111100101111101111001100111111001110000110110101100000001000101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6000

pattern = 30; // 6000
ALLPIS = 207'b110000110111000101110010101011100001001100000010010011000111000111001010000111000010110110010001101101101011101111100010011000100111110111010010101001101010000100101101101000001101101000101101011001000001010;
XPCT = 108'b110101000110110100010110101101000001110011110111111111011111000011011111001100010100111010111111111011000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6200

pattern = 31; // 6200
ALLPIS = 207'b011000011011100010111001010101110000100110000001001001100011100011100101000011100001011011001000110110110101110111110001001100010011111011101001010100110101000010010110110100000110110100010110101100100000101;
XPCT = 108'b001110100011011010001011010100100000100111111011111110011111100111011111011101011000110100011111100100001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6400

pattern = 32; // 6400
ALLPIS = 207'b101001100100100100100101100101100100101100010001101011011010001111111011100100100110010100110111110001110100000110100110101011001011100000110111101010011001100100110011011010000100010100100111111001010010100;
XPCT = 108'b111011010010001010010011111101010010110001110111110101000000101101100110011001000100101000111111111100111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6600

pattern = 33; // 6600
ALLPIS = 207'b000011111101101101101100111100111101100111010101110001101100101100000101011101101111110001111010001101101001000111001111000001111001011000111010010000111111111101111111101100100101010001101110000111000110001;
XPCT = 108'b001101101010101000110111000011000110010110111010001010011111111111011111111101010111110100011001101001010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6800

pattern = 34; // 6800
ALLPIS = 207'b101000011010010010010011111011111010011111111011010011101100011001111001001010010001101100001010110111000000100101000001001011110111001100101010100010000110011010001100101100010110111100010000111010110001100;
XPCT = 108'b110101100011011110001000011110110001101001111110100101101111100101010101111101110100110000000001001000011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7000

pattern = 35; // 7000
ALLPIS = 207'b011101101001101101101100011000011001100011101100000010101100000011000111000001101110100010110010101010010100010100000110001110110000000110100010111011011010101001110101001100001111001010101111100100001010010;
XPCT = 108'b000001100111100101010111110000001010110111111001111110011111101100101011000101110111111011100111010011011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7200

pattern = 36; // 7200
ALLPIS = 207'b101110110100110110110110001100001100110001110110000001010110000001100011100000110111010001011001010101001010001010000011000111011000000011010001011101101101010100111010100110000111100101010111110010000101001;
XPCT = 108'b111100110011110010101011111010000101000001111110001011010000101100011110010001001100100110111111110101100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7400

pattern = 37; // 7400
ALLPIS = 207'b101110001011001011011010001101011100000001011011000001100110011100001001000001101001001011110001000111000000010110011111011001000010011000100000011011010010010111011000111000010101101101000100111001010110100;
XPCT = 108'b110111000010110110100010011101010110001011111110001011111111100001111111110110110000110010011000010001101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7600

pattern = 38; // 7600
ALLPIS = 207'b010111000101100101101101000110101110000000101101100000110011001110000100100000110100100101111000100011100000001011001111101100100001001100010000001101101001001011101100011100001010110110100010011100101011010;
XPCT = 108'b000011100101011011010001001100101011000111111001011010011111100110111111110111100100110111000111000001100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7800

pattern = 39; // 7800
ALLPIS = 207'b001011100010110010110110100011010111000000010110110000011001100111000010010000011010010010111100010001110000000101100111110110010000100110001000000110110100100101110110001110000101011011010001001110010101101;
XPCT = 108'b001001110010101101101000100110010101000101111001011010001001001100001110100111110000111010000001101010101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8000

pattern = 40; // 8000
ALLPIS = 207'b101100010101111101111110110100001111001100011010110011010110111100011010101100101011011101101001111001001100000100010101010000000011110011110011101001000011110110001000011101000110111001001111011110011000010;
XPCT = 108'b110011100011011100100111101110011000100111111110101111111111110110000101111111100001111000100110100010100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8200

pattern = 41; // 8200
ALLPIS = 207'b111111101110011010011010111111100011001010011100110010110001010001110110110010110011111010000011001101010010000100101100000011001010011001001110011110111000011111110111010100100111001000000000010110011110101;
XPCT = 108'b111010101011100100000000001010011110010111111101011011100000111110010110000001011011101011111110100001000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8400

pattern = 42; // 8400
ALLPIS = 207'b011111110111001101001101011111110001100101001110011001011000101000111011011001011001111101000001100110101001000010010110000001100101001100100111001111011100001111111011101010010011100100000000001011001111010;
XPCT = 108'b001101010001110010000000000111001111011010111011011010011001111000001110100101000100110110000001100110110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8600

pattern = 43; // 8600
ALLPIS = 207'b000011001111100001000001100101001110001111011011010011111011001101110011000100000101010101001011100001010000010011110110110101111100100011010010000110111011110001100111010111100110110011010011111110011010100;
XPCT = 108'b001010111011011001101001111110011010010101111011010000001111111111111111011111110110111100011111100001010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8800

pattern = 44; // 8800
ALLPIS = 207'b001101100101001110100111001110000101011001101111101010001001111011011010100111110100001011111110110001011010000001001000010011110001011000011000111110111011101010110011000010111111110010000000111010011101011;
XPCT = 108'b001000011111111001000000011110011101111001111001111110011001100100100110000101001111111100100000101100001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9000

pattern = 45; // 9000
ALLPIS = 207'b000110110010100111010011100111000010101100110111110101000100111101101101010011111010000101111111011000101101000000100100001001111000101100001100011111011101110101011001100001011111111001000000011101001110101;
XPCT = 108'b000100000111111100100000001101001110011100111010001010001111011001011111101111111100110111000000100011011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9200

pattern = 46; // 9200
ALLPIS = 207'b000011011001010011101001110011100001010110011011111010100010011110110110101001111101000010111111101100010110100000010010000100111100010110000110001111101110111010101100110000101111111100100000001110100111010;
XPCT = 108'b000110001111111110010000000110100111000111111000000000011111100010111111010111100010110111111111001101011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9400

pattern = 47; // 9400
ALLPIS = 207'b100001101100101001110100111001110000101011001101111101010001001111011011010100111110100001011111110110001011010000001001000010011110001011000011000111110111011101010110011000010111111110010000000111010011101;
XPCT = 108'b111011000011111111001000000011010011101100111111111111000000101111011110010011111101100011111111011111111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9600

pattern = 48; // 9600
ALLPIS = 207'b010000110110010100111010011100111000010101100110111110101000100111101101101010011111010000101111111011000101101000000100100001001111000101100001100011111011101110101011001100001011111111001000000011101001110;
XPCT = 108'b001001100101111111100100000011101001110011111001111110010000100111111110000000100111100000011111100110100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9800

pattern = 49; // 9800
ALLPIS = 207'b000001111111101110111000101011111000100110100010110100001110011100001101010001101001111100100000001100010110110010100100111011101100000010000111011011100100010011100110111100000001101011000011111000100110011;
XPCT = 108'b001111100000110101100001111100100110100011101001111110011111001000101111001100011011110001100110110011111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10000

pattern = 50; // 10000
ALLPIS = 207'b001001011011010011111001110000011000111111000000110001011101000001111101001100010010101010100111110111111111011111110100110110111101100001110100000111101011101101000000000100000100100001000110000101000001101;
XPCT = 108'b000000100010010000100011000001000001100111111011110100001111010111011111011100000101110000111110100100010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10200

pattern = 51; // 10200
ALLPIS = 207'b101101001001001101011001011101101000110011110001110011110100101111000101000010101111000001100100001010001011101001011100110000010101010000001101101001101100010010010011011000000110000100000100111011110010010;
XPCT = 108'b111011000011000010000010011111110010110011111111111111011001100101001110001100010001111000011001010000111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10400

pattern = 52; // 10400
ALLPIS = 207'b010110100100100110101100101110110100011001111000111001111010010111100010100001010111100000110010000101000101110100101110011000001010101000000110110100110110001001001001101100000011000010000010011101111001001;
XPCT = 108'b000101100001100001000001001101111001010111111011011010001111010011100101000111000100111110100000100110000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10600

pattern = 53; // 10600
ALLPIS = 207'b000010110110110111110011110010111110100000101101110111100111000100001010110100001101100100101110110011010110111100110001100111001110110100110100110000000010100000010111101100000101110101100110110111101110000;
XPCT = 108'b001101100010111010110011011011101110010101101011011010011111010011111011001100100100110100000001010111110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10800

pattern = 54; // 10800
ALLPIS = 207'b100001011011011011111001111001011111010000010110111011110011100010000101011010000110110010010111011001101011011110011000110011100111011010011010011000000001010000001011110110000010111010110011011011110111000;
XPCT = 108'b111110110001011101011001101111110111110011111110101111011111110010011111010100100001110001011111001101011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11000

pattern = 55; // 11000
ALLPIS = 207'b011001001001001001011001011001001011000100011010110110100011111110111001001001100101001101111100011101000001101001101010110010111000001101111010100110011001001100110110100001000101001001111110010100101001000;
XPCT = 108'b001100000010100100111111001000101001100111111001111110011111110010100111100110110110110001111110001000101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11200

pattern = 56; // 11200
ALLPIS = 207'b001100100100100100101100101100100101100010001101011011010001111111011100100100110010100110111110001110100000110100110101011001011100000110111101010011001100100110011011010000100010100100111111001010010100100;
XPCT = 108'b001010001001010010011111100110010100110011111010101110010000110100111110100000011001100111111111110001101110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11400

pattern = 57; // 11400
ALLPIS = 207'b100110010010010010010110010110010010110001000110101101101000111111101110010010011001010011011111000111010000011010011010101100101110000011011110101001100110010011001101101000010001010010011111100101001010010;
XPCT = 108'b110101000000101001001111110001001010011101111110001011011001001101111110000101000100111101000000011110010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11600

pattern = 58; // 11600
ALLPIS = 207'b010011001001001001001011001011001001011000100011010110110100011111110111001001001100101001101111100011101000001101001101010110010111000001101111010100110011001001100110110100001000101001001111110010100101001;
XPCT = 108'b001110100100010100100111111010100101000011111001011010011111110011001111110110110000111111011111111001010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11800

pattern = 59; // 11800
ALLPIS = 207'b010001000100100100111001011101101001010000110010101010001000010101010010111011011111011000010100101000100111110110111110000110010000000100000101010101011001011110010011100011111111101000011100010001011101101;
XPCT = 108'b001100011111110100001110001001011101111010101001111110000110000011011111111011111110100111111111010100111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12000

pattern = 60; // 12000
ALLPIS = 207'b101010101011011011101110010101100110001001111100000001010100100000001100101011010001011100100011000101011100010110100011001111101000001010001000000000011110010011101110110110000000100100110110101010010101100;
XPCT = 108'b111110110000010010011011010110010101000011110110001011101111101010101111011111011000110110111111110111001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12200

pattern = 61; // 12200
ALLPIS = 207'b010111011100100100000101110001100001100101011011010100111010111010100011100011010110011110111000110011100001100110101101101011010100001101001110101010111101110101010000011100111111000010100011110111110001100;
XPCT = 108'b000011101111100001010001111011110001001111111001011010000000010010001110101001101000101100111111010000100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12400

pattern = 62; // 12400
ALLPIS = 207'b101001100111011011110000000011100010010011001000111110001101110111110100000111010101111111110101001000111111011110101010111001001010001110101101111111101100000110001111001001100000110001101001011001000011100;
XPCT = 108'b111001001000011000110100101101000011110001110100100101101111000101101111110101000001111010011111101101111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12600

pattern = 63; // 12600
ALLPIS = 207'b010100110011101101111000000001110001001001100100011111000110111011111010000011101010111111111010100100011111101111010101011100100101000111010110111111110110000011000111100100110000011000110100101100100001110;
XPCT = 108'b001100101000001100011010010100100001111111111011111110011111001101110101100110111100111001011001011010110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12800

pattern = 64; // 12800
ALLPIS = 207'b000100001000011111100111011101110101000010101011101101111001111011101100011011100101110111101010000001100000001101001011010001011001010101110000111010100100111110100010011010110011101110010001011010010101110;
XPCT = 108'b001011011001110111001000101110010101101001111011111110000000111100000100111000000001100010111000100001010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13000

pattern = 65; // 13000
ALLPIS = 207'b010000000110100011000000101010110100000000011000010001010110001011101001111101100110000101101110001000111111110101101100110010000110010001011001011011110000010001111011000101010011010011111000000111111000110;
XPCT = 108'b001000100001101001111100000011111000111110101011111110000000100100101010000000101101101101111110110000110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13200

pattern = 66; // 13200
ALLPIS = 207'b000110001000100001000010110001111111100001100011010000000101001000011111101001100111010001110010110011000000010000100111000000000001101100011100111100001110111000111001110110101011100100000110100011000101011;
XPCT = 108'b000110111101110010000011010011000101010001111000001010000000100110101110001000101010100110100110010111000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13400

pattern = 67; // 13400
ALLPIS = 207'b100001001101011001010011100011101101010001010100111100010010001110101010000010001101011000010000001000101111100101101111101100100000111110000100110100110101100000111011111100101010100010111011110011011001111;
XPCT = 108'b111111101101010001011101111011011001110001111100101111101001100101101110100101111011110111100111000100101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13600

pattern = 68; // 13600
ALLPIS = 207'b111010011010011111100110000011101001110101110000011011010100001001001111010110011101100110101101010011000100010100100111110111101000000111101011100111111111100100101001111000110101111000010110011110001101001;
XPCT = 108'b110111001010111100001011001110001101011111111111011011011111000010000101100101000000111000000001101001001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13800

pattern = 69; // 13800
ALLPIS = 207'b111101001101001111110011000001110100111010111000001101101010000100100111101011001110110011010110101001100010001010010011111011110100000011110101110011111111110010010100111100011010111100001011001111000110100;
XPCT = 108'b110111100101011110000101100111000110101111111111111111001111111010111111011100010000110001111001111000011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14000

pattern = 70; // 14000
ALLPIS = 207'b111100101111101110001011011011101000111100111001010010100101101000110110000011011001101001000010000101111110101000110101110001011010001001110000010011001101000101101101011001110010001110111101000101011000000;
XPCT = 108'b110011001001000111011110100001011000111111111101111111101111111011011111101111000011110011011000011111000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14200

pattern = 71; // 14200
ALLPIS = 207'b111100011110111110110111010110100110111111111001111101000010011110111110110111010010000100001000010011110000111001100110110100001101001100110010100011010100011110010001101011000110010111100110000000010111010;
XPCT = 108'b110101010011001011110011000000010111110011111111111111010000100111001110001011110100100101100110111100111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14400

pattern = 72; // 14400
ALLPIS = 207'b111111000111101111101101110101101001101111111110011111010000100111101111101101110100100001000010000100111100001110011001101101000011010011001100101000110101000111100100011010110001100101111001100000000101110;
XPCT = 108'b110011011000110010111100110000000101001011011111011011001111000011101111110110110001110110000001000100011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14600

pattern = 73; // 14600
ALLPIS = 207'b011111100011110111110110111010110100110111111111001111101000010011110111110110111010010000100001000010011110000111001100110110100001101001100110010100011010100011110010001101011000110010111100110000000010111;
XPCT = 108'b001001100100011001011110011000000010001011111011011010001111010011011111111100000101111101100110011010111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14800

pattern = 74; // 14800
ALLPIS = 207'b110101110001110100001111010101111111101100011010100111101010101110011000001011010000010100100001000001101000001100001111000001001000010010010011001111110100010100011011100100101001011100010111101110111011111;
XPCT = 108'b111100101100101110001011110110111011110111111111111111001111101010011111000101110101111110011000001111110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15000

pattern = 75; // 15000
ALLPIS = 207'b011000110001110011110101010001101101010111101000000111100101111101101001110011010110111010111001110001111011101011111011101100000100000001000011001101001000110110101010110101101011111110110011010101100110101;
XPCT = 108'b001110101101111111011001101001100110100111111011111110011111101100101111111100011000110000011111110000111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15200

pattern = 76; // 15200
ALLPIS = 207'b000111001000111000000100001001110010000101001000101011110001001010001000100111101010110110111010110100111001001100000000111101010001000100010101100110001011010011111001001110100101010111110000100100000100000;
XPCT = 108'b000001111010101011111000010000000100010101111010001010010000111110001110010000000110100100111110101010000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15400

pattern = 77; // 15400
ALLPIS = 207'b000001101101010101110000111111101011100011000001000001101000001111100001100101001011101011110100001011010011001011111100010010001000101010000000011001110111010101011011100000101101111011000000110000111001010;
XPCT = 108'b001100001110111101100000011000111001110001111010101110011111010000011111111111110100111100011111101011101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15600

pattern = 78; // 15600
ALLPIS = 207'b000000110110101010111000011111110101110001100000100000110100000111110000110010100101110101111010000101101001100101111110001001000100010101000000001100111011101010101101110000010110111101100000011000011100101;
XPCT = 108'b000110000011011110110000001100011100111011111000100100001111010111111111001100101010110000100001111011101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15800

pattern = 79; // 15800
ALLPIS = 207'b000100010010010011100101110110100101000011001010101000100001010101001011101101111101100001010010100010011111011011111000011001000000010000010101010101100101111001001110001111111110100001110001000101110110101;
XPCT = 108'b001001111111010000111000100001110110101101011000101110011111111000101111110101100111111110000000011101011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16000

pattern = 80; // 16000
ALLPIS = 207'b010000010001111010101101101101111110011101111001000010011101101100001101111001110110101111100101000101010110100010010111100110001000011110111111000101010010010001010111000000010000100111101101010000110100000;
XPCT = 108'b001000000000010011110110101000110100111011111001111110011111110010011111001111111111110110111111111010111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16200

pattern = 81; // 16200
ALLPIS = 207'b110010111000111101110101101101010010011011011000101111111011101111110001011001101110010010100001000101111010000011100001100101101101101111101001010101110101101001011000011000111011111111111100110011000000100;
XPCT = 108'b110011001101111111111110011011000000001011111111011011001111000000111111101111000001111111000001010110000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16400

pattern = 82; // 16400
ALLPIS = 207'b101100001101111010000110000000101000011101000100001111000101100011100111100101110110111011100010011011110011100100010111010101001011100110000100011111111001111000111000000110101111110000100101101101011000001;
XPCT = 108'b110000111111111000010010110101011000100101111110101111101111000001011111110101001101111100111001110000010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16600

pattern = 83; // 16600
ALLPIS = 207'b111011100000101011111010111011110110111100100011000111001010000000100010001010110000110001110010101100010001111101101010111001000010000100011111001101011010111100100000000001001010110011010011111010111110000;
XPCT = 108'b110000000101011001101001111110111110000011111111011011010110100111001111100010111111100111011110000010101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16800

pattern = 84; // 16800
ALLPIS = 207'b001111111111110000000100001100100010001100010110011100000010001000011111100010111011011001000100011111001111001011000010011011011000101101011101110011001111110101001010000000101000011001000000111110111111110;
XPCT = 108'b001000001100001100100000011110111111000101111000001010001001010100111110110100011111111010011000110011111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17000

pattern = 85; // 17000
ALLPIS = 207'b100011101110000110101100101110110110111110111100100101011101001110001010000001011000011001110100000010100101010000100111000000111110010101101000011001100001101100000101100000011010100001111101011111011011111;
XPCT = 108'b110100000101010000111110101111011011011111111111011011101001110110111110010100100010110100100001101001111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17200

pattern = 86; // 17200
ALLPIS = 207'b101000101010011011000110100110010011110010010110001011001010111111101111011001100000101001111000000101111111110110011110010110000111111011100101000011001010001010010110011000010110001111110010000111000010111;
XPCT = 108'b111011000011000111111001000011000010101101101111111111111001100101101110010110000001110011000001010110101001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17400

pattern = 87; // 17400
ALLPIS = 207'b010111010111000101001000111011111100110011010101110100100010100011011101101111100000011111010110001001110100100011011011111001111111001011101111000011111000100010001011100100110110100001011001011010000101100;
XPCT = 108'b001100101011010000101100101110000101011011111001011010001111110001111111011110101100111100011110010001010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17600

pattern = 88; // 17600
ALLPIS = 207'b010000111101000111011011001001100100001110100110010100011010111101001110010001110101011011010001000011111000011110111000010000111111000100111001000111011000010010011100010001100101110011100101110111010001110;
XPCT = 108'b000010001010111001110010111011010001100111111001111110011111110111101111011100111011111100111111010010111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17800

pattern = 89; // 17800
ALLPIS = 207'b000100011110101011011011011111100111011110010000100111011011000011011110011101101011111001010001010101101000100101111001100010000111101111110001010100100100010101110000000100001001111011010100001101000000011;
XPCT = 108'b000000100100111101101010000101000000100111111011111110010000000010111010011001001101101000111110101101111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18000

pattern = 90; // 18000
ALLPIS = 207'b000001000111101010110110110111111001110111100100001001110110110000110111100111011010111110010100010101011010001001011110011000100001111011111100010101001001000101011100000001000010011110110101000011010000000;
XPCT = 108'b000000000001001111011010100011010000100001111010100100011111100100011111001101101101111111111111010000010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18200

pattern = 91; // 18200
ALLPIS = 207'b011101000000100011010101010111011100000000011111111000011111111101110111101000111001001010110001110011010000001000100100110001000001001011111000001000100011110100000010011001110111001101011000000001111110110;
XPCT = 108'b001011001011100110101100000001111110101011111001111110000000111011101110110000100011100011111111010100010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18400

pattern = 92; // 18400
ALLPIS = 207'b010101000100111000000111111100011000110000010110000101110110000011100110111000001000011001101110010001000001001110011101110110110101111000010101101110011000111100010011111010110110000100010111100001011001111;
XPCT = 108'b001111011011000010001011110001011001111010111011111110000000001011001110111000010001101000100110011110100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18600

pattern = 93; // 18600
ALLPIS = 207'b001011000100111000000000011101011010100011011001011110001111011010100100001001010111111001111011010110100000001110010100001010001010001110100111011100010010101010110011110000000001100110011111011111100100111;
XPCT = 108'b001110000000110011001111101111100100010101110001011010001001110011101110101111110100111011000000100101110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18800

pattern = 94; // 18800
ALLPIS = 207'b101001100110010000101111111110100011110101001110110000110100011111010011000110000000011000000111010011110001000110000111111100100100100011011111001000100001100010010100001101000110010110110110111110011111111;
XPCT = 108'b110001100011001011011011011110011111100111110101111111100000011110001110100010010101101101111111110110011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19000

pattern = 95; // 19000
ALLPIS = 207'b110100111001110101100001010100000110111101011100010000000010111001001111000101111100100011011001001101010100010101110011100111101001101101001011110110011001100010100100001111101010000011000001101111011000100;
XPCT = 108'b110001111101000001100000110111011000100111111101111111001111011110111111011110100111111111111111010001011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19200

pattern = 96; // 19200
ALLPIS = 207'b100111011100011001100101111101011111011110110001110000011110100001010000001010000111011011011101010101111010000010011101000010110101111101011101110011101111000101010000011110000010001100111000110110010010100;
XPCT = 108'b110011110001000110011100011010010010000101111101011011100000111011110110101000111001101100111111001001001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19400

pattern = 97; // 19400
ALLPIS = 207'b110111010111010111110011110100111001110111100011100000001000010110101111110110111101010011101111101100110110100100110101001000001101111010101011011000101010001011010101001011011011000101100010001101011011110;
XPCT = 108'b110001010101100010110001000101011011011111110101011011001111101001111011000111110010110010000111110111101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19600

pattern = 98; // 19600
ALLPIS = 207'b011011101011101011111001111010011100111011110001110000000100001011010111111011011110101001110111110110011011010010011010100100000110111101010101101100010101000101101010100101101101100010110001000110101101111;
XPCT = 108'b001100101110110001011000100010101101000111111001011010001111001000101111010100110100111100111000110101110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19800

pattern = 99; // 19800
ALLPIS = 207'b101101110101110101111100111101001110011101111000111000000010000101101011111101101111010100111011111011001101101001001101010010000011011110101010110110001010100010110101010010110110110001011000100011010110111;
XPCT = 108'b110010011011011000101100010011010110111011111101111111001111110001011111000100011011111101100001011010010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20000

pattern = 100; // 20000
ALLPIS = 207'b010110011101111110001010011000001111100111000001110110011111011100101101010111100010111111111111001101100011010010110111100101100001111100010010100101000001011100101111001101011010100001001110001001001011011;
XPCT = 108'b001001100101010000100111000101001011011011111001011010011111111010101011000110010111111110111001100100101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20200

pattern = 101; // 20200
ALLPIS = 207'b110110001110011100010000011011011011110011111111000011010000010011100001000011001000010101001110010101100001100001111111000011110001110101110001011010000011011010010101111111011010011101111111000101011011011;
XPCT = 108'b110111110101001110111111100001011011011111111111011011000110100111111111101001000000100001100111101000100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20400

pattern = 102; // 20400
ALLPIS = 207'b010011000011110110101110101101011000111100110000001100111011111010000011100100101110100000001011011100110000011100001101101000011100111000100000010010110001001100100100010011001101000001110011110001101001101;
XPCT = 108'b000010010110100000111001111001101001000011111001011010001111100101011111110100101110110010111001011011100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20600

pattern = 103; // 20600
ALLPIS = 207'b010000001000110101010101110111000000000111111110000111111111011101111010001110010010101100011100110100000010001001001100010000010010111110000010001000111101000000100110011101110011010110000000011111101100010;
XPCT = 108'b001011101001101011000000001111101100101111111011111110000110100101011111111011110001100100011111101100011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20800

pattern = 104; // 20800
ALLPIS = 207'b101010010000010110010001011110011101001011110000110001001011000010010100001101111011010011100111101000111010000000000011011000111111110110100010111111100101010010000010111010011000001111100010100110110010100;
XPCT = 108'b111111010100000111110001010010110010001101111111011011011111000011011111010101110000110011000000100111100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21000

pattern = 105; // 21000
ALLPIS = 207'b110101111011111111110101000111011000011110010010100000101110100100100000100011000000100011100110111000110101111101010110011100001111000100010111011000101011100101110101011101100111000100010011000011101110000;
XPCT = 108'b110011101011100010001001100011101110110011111101111111011111001010111111010100100100110011011000001011000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21200

pattern = 106; // 21200
ALLPIS = 207'b010101001011111000010110110110010010001110001110111100000010111110100111111001010011100001000000011011101111110101111100101101011010011100111000010000001110101110100000110101101100101000111001001000000110011;
XPCT = 108'b000110101110010100011100100100000110100011101001111110011111011010001111001100001110110000100110000101111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21400

pattern = 107; // 21400
ALLPIS = 207'b110101010010111110000101101101100100100011100011101111000000101111101001111110010100111000010000000110111011111101011111001011010110100111001110000100000011101011101000001101011011001010001110010010000001100;
XPCT = 108'b110001100101100101000111001010000001101011111111111111101001111101001100010101110010110100100000011000011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21600

pattern = 108; // 21600
ALLPIS = 207'b000001111111101101011010011011011010011001001100100001110011100110100101011001111001110111010110000001110001001000010100111001011110101011100100101100001111011001111000100110101100010110000001110101010010010;
XPCT = 108'b000100111110001011000000111001010010100111111010101110011111100011110111000101101011111101000000001111000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21800

pattern = 109; // 21800
ALLPIS = 207'b111000001101100101000100111011111010001010101110011011110111001101000010101000001001101111010110000010000101010010001111110100100101001111011011110100000101101011010010111001110010000111100101001101101100100;
XPCT = 108'b111111001001000011110010100101101100101111111111111111101111000000111011011101000000110111111110000101110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22000

pattern = 110; // 22000
ALLPIS = 207'b000010101000111101011100111100100001001101010010100001001010111101111110001100011101001111001110101100010101010101001001010011001101101111101100110000100010111111101100010110101011001111101111000111101111100;
XPCT = 108'b000010111101100111110111100011101111000111111010000000001111100000011111111111111001110010000000101010110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22200

pattern = 111; // 22200
ALLPIS = 207'b100011110010111111110110110011100111111011101011001110010000001101011000100011111111110110000010101000000011101011000100101100101011011010111010111000101110110000010000100100110001000011100100010011101001011;
XPCT = 108'b110100101000100001110010001011101001001001111101011011010000011000101110101001101010101111111110001001001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22400

pattern = 112; // 22400
ALLPIS = 207'b110001111001011111111011011001110011111101110101100111001000000110101100010001111111111011000001010100000001110101100010010110010101101101011101011100010111011000001000010010011000100001110010001001110100101;
XPCT = 108'b110010010100010000111001000101110100101011111111111111101111010111001111111111011111110110111001110001011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22600

pattern = 113; // 22600
ALLPIS = 207'b010100111000000100001111011101100011100111001010110110000101001000010111011000110000001111111011011100100010101010111011100011000110101100100010100001010000111111011101111101110110110110100001001111101001000;
XPCT = 108'b000111101011011011010000100111101001111111111001111110011111110101101111101101000010110100100001110001000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22800

pattern = 114; // 22800
ALLPIS = 207'b101110011101110000011011100010101000001011001101010110101100011010101111110110100011001011011101101111110001011011011110001001101101110110100110011100100000011111101001011010001010001000000111010011101101101;
XPCT = 108'b110011010101000100000011101011101101010011111100001011111111001111111011000100100011111100011001111011000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23000

pattern = 115; // 23000
ALLPIS = 207'b110111001110111000001101110001010100000101100110101011010110001101010111111011010001100101101110110111111000101101101111000100110110111011010011001110010000001111110100101101000101000100000011101001110110110;
XPCT = 108'b110101100010100010000001110101110110000011111111011011000110111110011101111001110010100100111111111010101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23200

pattern = 116; // 23200
ALLPIS = 207'b111110000001010001110101101111110010111010110010100100100101101110001101011101001011101111011001000101111101100000011111011101100110110100001110001011001010110011101101101111100000010010100100101001110100110;
XPCT = 108'b110101111000001001010010010101110100010011111101011011100110011110011111000001110110101110011110110010111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23400

pattern = 117; // 23400
ALLPIS = 207'b010101100010110001001101110100010000000000010000111001010001001000111110101100101000010100011111000011010101011111100100100000100101111101110011000100100000011000100100100111111010100110100001111101010000111;
XPCT = 108'b000100111101010011010000111101010000101111111011111110000110011100111111001000110100101001000111001101111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23600

pattern = 118; // 23600
ALLPIS = 207'b111101110100001001101000101001100100000101100010101001001101101101000001110000001001011010100010100011100101101000111110011001110111010001010011001100001011010001100110100010000111101010000010100111111010000;
XPCT = 108'b111100010011110101000001010011111010100111111111111111110000000010001110010000111100101010111111100011010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23800

pattern = 119; // 23800
ALLPIS = 207'b111111100001010000110011101110001101100001111100011100111000000110001101110000111111101101011011100111111000110110010001001100111111111110000000110000001010000101010111001110111100110001011100001001100001100;
XPCT = 108'b111001111110011000101110000101100001011011111101011011101111011101111101001100110111111101011001010101001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24000

pattern = 120; // 24000
ALLPIS = 207'b011111011011100101011000001001110101111010011011100010000110001011110101001101001111001100111010010001110111010111010111000110001111111101100001011100011100101110101100100000101010011111110011011000111010111;
XPCT = 108'b000100001101001111111001101100111010000011111001011010001111101101111111011100101110110010111001111111110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24200

pattern = 121; // 24200
ALLPIS = 207'b111011001001010101010101101010010011011100010101101011111100111110000011110000001001010101111101101110000011001101010000000111010001111100101101110011110010101101110000011110100010101001101000001100110100100;
XPCT = 108'b110011111001010100110100000100110100000110111111011011001111100010101111001101010100111011011000111010001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24400

pattern = 122; // 24400
ALLPIS = 207'b100001110000110100110010000110111111110100111101100011001111000011111011011101111101001111101000010100010001011111110110011000001011100011001010111100101000100001110010011010010001001000100010010000001110001;
XPCT = 108'b111011010000100100010001001000001110101001111111110101110000111110001010011001011110100011011111100010011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24600

pattern = 123; // 24600
ALLPIS = 207'b111011101101101011001111000001100000011000001000010011001000000000100110011111101101101000101111001101011001011001111010010111100101101111001110010001111010111101111101110111000111110001110111010101000111011;
XPCT = 108'b110110110011111000111011101001000111010110111111011011111111000100001111000111110101111010000001111101011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24800

pattern = 124; // 24800
ALLPIS = 207'b000110100100000010011011011011010011010010001010111011110010011001010001100101100000011010010000000101101111110011001000000111110000110110011111010100111000111000101001001111110101000100101001110000111000011;
XPCT = 108'b000001111010100010010100111000111000011011101010001010010000011000111010001000000101100111000111011100000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25000

pattern = 125; // 25000
ALLPIS = 207'b110111011100001000010001101000100001111101101011100011111000010110100011000000001110011010011001010111111010011010011001001010111101111101111110101111010111000100111011110000000001000011011010111101111001000;
XPCT = 108'b111110000000100001101101011101111001010111111111011011111001110111101010000101100000110000100000000000111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25200

pattern = 126; // 25200
ALLPIS = 207'b011001111100101010101011011100011110011000101010001110111110011010100001101100100101010001111011001101101010101000100111110100101000110000000110001010000011010100011101000011111110000101010000101000110111001;
XPCT = 108'b000000011111000010101000010100110111111011111001111110010110000110011111110011011111101001011111110100110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25400

pattern = 127; // 25400
ALLPIS = 207'b010111011010011101111100010110010101011010010100011110011000000110101101100011100101011011001100010101101000010011011000100000010011011110111001101011110101110000100010111011100010001010001100001000101111101;
XPCT = 108'b001111011001000101000110000100101111000011111001011010000000010001101110100000001110101010111110111011100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25600

pattern = 128; // 25600
ALLPIS = 207'b100101111101111001010101011111111100001110110100011111111111100101000011100100011010110001000110000110001000001011010111010110111001010010000100010001110111111100100000010010101110110111100010010011010011111;
XPCT = 108'b110010011111011011110001001011010011100001011111111111001111101101101011111100100001110110000110110010010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25800

pattern = 129; // 25800
ALLPIS = 207'b011010011010100100101110101111110111110101111101111110100011101100100000011100011001110001011111011100111110111101101110101110011101110101110110001101010111110000010011100010110001111110110011111010010111110;
XPCT = 108'b001100011000111111011001111110010111011011000001011010010000100011011110011011111101101111111001101111010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26000

pattern = 130; // 26000
ALLPIS = 207'b110011100010100001010101100001101011111001000011111000001111010101001001010100000011101111000101111010000011111110011001111101110010110010000100111010111011011011001111001010101011010000100100111101001100110;
XPCT = 108'b111001011101101000010010011101001100010111111101011011100000001000011110011001101111101101100110111000001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26200

pattern = 131; // 26200
ALLPIS = 207'b110001001010000011000100010011101110100101101110001011100110011011110110110000000001001010111010101111010110011110001111100111000111111101000001110111100110110010100010101111010100100010111010001100110001100;
XPCT = 108'b111101110010010001011101000100110001101111111111111111100000101110011110001011101001101110111111010111011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26400

pattern = 132; // 26400
ALLPIS = 207'b111000101011001101111001011000101001100001000000101100010110101010011000001110000110011110101110101110111010000100001010101111110111101110101001001100001011000001110100000110110010101100111101110000111111110;
XPCT = 108'b110000111001010110011110111000111111101011111101111111101111011010111111010101111111110010100000000011010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26600

pattern = 133; // 26600
ALLPIS = 207'b100111110101100011100011001001101011101000100011100110000011100010100011100111100010001101111110100000110111011010111011110010101110110111100001100011010110111001001101110110110111100101011100010011010000110;
XPCT = 108'b110110111011110010101110001011010000011001111100001011101111101100101011101100111001110100000001000010111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26800

pattern = 134; // 26800
ALLPIS = 207'b111101101110000001001010101010100011100101001110110001011100010011110001101111010111110111111000100001101000011111011101111010010110000010000011111111101110101010110101111110111110100011101111010111100001101;
XPCT = 108'b110111111111010001110111101011100001111111111111111111000000110111101110001000000000101111011110111011111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27000

pattern = 135; // 27000
ALLPIS = 207'b110101101011110001110110011101011011110111110001011010100101000100110100011111000001011010100001101110010101000011001010000010011101010001010110000100101010101100001011011101110110101110011101110101010011111;
XPCT = 108'b111011101011010111001110111001010011111111111101111111101111111010111011100110101000111110000111001101111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27200

pattern = 136; // 27200
ALLPIS = 207'b010100011011011100111000011011010011000010010001111010010101001111000111000100111010010001111000110100111011111110110110100011001100110110000000011101100101001110110111011100101101110011011101010001001111100;
XPCT = 108'b001011101110111001101110101001001111110011111001111110011111110011001111101111110011111011111111100111011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27400

pattern = 137; // 27400
ALLPIS = 207'b001001100010110011010100011011101011101110000110001101100100110111000000101111011000011011001100011011100011110000101011010110000110011010100011111110101010100100011011001010001000001010010001101101010100110;
XPCT = 108'b001001010100000101001000110101010100110101111010101110000000001001001110111001111111101001100110011110111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27600

pattern = 138; // 27600
ALLPIS = 207'b000100000100110111011100111000010001010010010000100010000001101011111100000100001110011100011110011010010101111111111000011101010011100001101101111000000010111101111010110101011001111110111000010101101111001;
XPCT = 108'b001110100100111111011100001001101111101111111000100100001111000110111111011100111010110000000001101011010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27800

pattern = 139; // 27800
ALLPIS = 207'b100011000010010100110001001101000010011111100001111001000000110101001101110011011001011000001111010111110101000001000010010000000000100100011001100110000010111001011110100110111101111110011110110100001011101;
XPCT = 108'b111100111110111111001111011000001011001101111110001011100000101111010110000011011110101101111110101100110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28000

pattern = 140; // 28000
ALLPIS = 207'b011001000100110111110101101000011001100011100000111000101001010000010110101111011101110101100110110110011110011010110000010010111011101110101010111110111100111100101101011011111011101100011101010000010010110;
XPCT = 108'b000011011101110110001110101000010010111011111001111110000000111010001110001000001110100000000110110011111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28200

pattern = 141; // 28200
ALLPIS = 207'b000111001111101110010100101100011010011011111001111000100000000010100101011110001110010001010001000011111000001000010110100010011000100101010011010000011100010011000000100101000001000010001111100001111100100;
XPCT = 108'b000100100000100001000111110001111100000001111001011010001111011110011111110101100100111000111110001100111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28400

pattern = 142; // 28400
ALLPIS = 207'b100000010101010101110100011110011000001110110010111101011000100101110011111000110111100001011101101101011101101010010011001011110110100111010110000011010001110110000000001010100011000010100100100010011101001;
XPCT = 108'b110001011001100001010010010010011101100001111111110101011111100010001111010111100101111110011111010101010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28600

pattern = 143; // 28600
ALLPIS = 207'b010000000111001010101010101011111101000000101101101000001101111100000000111101010011110010010111111010111110110111011100110011100101010011111110001000110111010001010111100111010011001010000000111110111101101;
XPCT = 108'b001100110001100101000000011110111101111111001001111110001111000010001111100110111110111010111111111111110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28800

pattern = 144; // 28800
ALLPIS = 207'b101001110010101101110100010001000001101000100011010111010011010011001001000010101010010011110000101110110000001110001010101010001101110111000010101101011110010011010110111101111011111100000001101010100110111;
XPCT = 108'b111111101101111110000000110110100110101001111111111111000000001100111110101011001101101010011001000010001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29000

pattern = 145; // 29000
ALLPIS = 207'b110001100010100111110111011001000100000000011101010110001010100000101111101100100010001001000101101011100100010100010100111011111011001011111000100101100100001110010000100100010001001010111000001010001101101;
XPCT = 108'b110100100000100101011100000110001101101011111101111111101111011100000111110110011101111101100000100011111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29200

pattern = 146; // 29200
ALLPIS = 207'b101000010000110110000111011100001111011101110011001111110001011000001101011110011011101100101110011110100101101101100110000111100011101011111101111100011010100010001001111001011011010101101010101000100011010;
XPCT = 108'b110111000101101010110101010100100011111001111110101111111001010000111110001100010000110101100000001100001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29400

pattern = 147; // 29400
ALLPIS = 207'b100000101010110010110011111000011001000000101010001110111000111100100110010100110110000001101110111011011110111110100010110111010101001110101101000100101001011101100100100000101010110101000000111001101100010;
XPCT = 108'b110100001101011010100000011101101100100001101101111111011001110000000100110100111110110100100001111110111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29600

pattern = 148; // 29600
ALLPIS = 207'b010111001110010110101111111100000000001010001101100111000011110101100011101000010011001111110100111011111110001011111000000111111101000011110001101011101010001100111100111001110110011000111000110000111011101;
XPCT = 108'b000111001011001100011100011000111011001011111011011010000000010111001110111011001111101010111111110100000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29800

pattern = 149; // 29800
ALLPIS = 207'b111011011010101011011111111001110000000100010111110011101001111111011001000110111100110011011000000111100101011000001110110001011010100100010100111110100011010001101001101100100111010101001100001110110010100;
XPCT = 108'b110101101011101010100110000110110010010111111111011011000000010111001110100011010110100000111110000111111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30000

pattern = 150; // 30000
ALLPIS = 207'b011101001110001100100011100110110111100010110010111011001101011011000010010011000011000110101101101000100101111011101100011100101111000010111001001111101101111011101110110011001100000000000101001010100101001;
XPCT = 108'b001110010110000000000010100110100101100011111011111110010000001001011110111011111000101111111111010101001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30200

pattern = 151; // 30200
ALLPIS = 207'b000011001110101100101110101010010111000111001001111111010001111001111111001100001100100000111001110001010001011010011010100011001011111100100110011000000110011101101100110110001101010101111100001101011001101;
XPCT = 108'b000110110110101010111110000101011001000111011010000000000110111010001111001000011011100110111111101111100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30400

pattern = 152; // 30400
ALLPIS = 207'b001011101101111011110100111010110110000010011001100001101100000111100110011101101001011101001010101111011110010110101001110001100010111011001011010001010010110100010011011111111001110010001011011000101100000;
XPCT = 108'b001011111100111001000101101100101100011001111011011010011111111111111111001100001110110011011001101100111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30600

pattern = 153; // 30600
ALLPIS = 207'b010101000101000011011100101110111110011010100011010001010100111101101000010010110011111000110001010001010100011010101101101001101101000101101110001001110010010011101101110011111110001111000000110101110101100;
XPCT = 108'b000110011111000111100000011001110101111111111011111110001111001111011111000110111110111110111001010110111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30800

pattern = 154; // 30800
ALLPIS = 207'b011000101001100100100101110001101011001100111011011000110000001001011111100011110010000001111100000001110010010001000100011001001001001011001111011000111100110011001000011110000000101101101010000110000010100;
XPCT = 108'b000011110000010110110101000010000010100111111001111110001111000000001111111111110011110010111110101100010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31000

pattern = 155; // 31000
ALLPIS = 207'b100001000111111110010101010111001101010100110100001001001110110101000100101000000111010010011100011101101100010100000000010000110111001111011110011010010000100001101011100100001100111101111100100110100100111;
XPCT = 108'b111100100110011110111110010010100100110101111110101111001001001011011110100101001001110001111000100011100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31200

pattern = 156; // 31200
ALLPIS = 207'b001010011110110010011001100000001100011000010100101110000011111000100010001000001110001110111010111010000111011000001100010001011001100001011110100000000000101101011111101001000001111111010110110100111011101;
XPCT = 108'b001101000000111111101011011000111011010111111000001010001111000110111111110111110101111111100001000010100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31400

pattern = 157; // 31400
ALLPIS = 207'b010101001000100000110011001010111011101010000011001011100100000101111110000000101011001101010000001111001011011011101000011110010000111110111001000111110111011101100101110100000111010001101000010000110111001;
XPCT = 108'b000110100011101000110100001000110111110011111011111110011111011101011111110111000011111111100001011010100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31600

pattern = 158; // 31600
ALLPIS = 207'b000001100111011111001001000000010001111010001110101100101100100100011010011110001011101010000000001011000101100111101010100110011110101101110000010001011010010010011011101101010000100011010010100001010111111;
XPCT = 108'b001101100000010001101001010001010111111010111000101110001111000001001111101110101110110111000110111001011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31800

pattern = 159; // 31800
ALLPIS = 207'b100001101110011101001011001111001000110011011010101001010010011111011110110010000100100011110000101101011101100010111001011100011101101101101010101000000101110000001001011111101101110010111011100001101110100;
XPCT = 108'b110011111110111001011101110001101110110011111110101111000110100111111111001010011000100100011110010001100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32000

pattern = 160; // 32000
ALLPIS = 207'b010001110100100010001110110011010000111001100000111111000010111100010111000001000110111011011001011110101001100100101001011100011111010100100011110001101101101111111001101111100110111010111011101110001011100;
XPCT = 108'b000101111011011101011101110110001011110111110011111110000110100011111111000000000110101101011111111000101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32200

pattern = 161; // 32200
ALLPIS = 207'b011001000001101111111110011101010100011011000000100001010100010100100101101110011101011111111101100111110010111110001100001011011010001100000010011011111000110010001000011100001011000111101101011100110001011;
XPCT = 108'b000011100101100011110110101100110001100111110011111110011111010010001111100100000010110001000111110000011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32400

pattern = 162; // 32400
ALLPIS = 207'b011010100010000101101001010110110001100101001100110111010111111101010001101011011110010010110100111111000010011110001001000101001111101111011101100101001011101000110010001011001101101110000101111100010111010;
XPCT = 108'b001001010110110111000010111100010111000111111011011010010000001111111110010011110101100001111001101011001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32600

pattern = 163; // 32600
ALLPIS = 207'b111111010010000101111011000000111110011100110011010100111011101110011110011110100101101101110111101011101100010101111011100000011110110110000001111101011010100101011010000100001010010000010101100010011001101;
XPCT = 108'b111000100101001000001010110010011001000011111101011011100000101100111110010000001111101110011110100111000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32800

pattern = 164; // 32800
ALLPIS = 207'b001110111001101010111001101100100011101010011111010110111111011111110001110010111011100110101110100111100111001101111001110011010101110011011000000111001001011101011000100110100011101110110011000000010011110;
XPCT = 108'b000100111001110111011001100000010011000011111000000000010110110011001111010001101110100010111110110010001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33000

pattern = 165; // 33000
ALLPIS = 207'b010111000010011111100001010010011011100100001001011011101011110000000110010010000010111000011100000011000100000011010101101100110111011101011110111100000111000111010111000111111001011100111111101010001110100;
XPCT = 108'b001000111100101110011111110110001110011011111011011010001111100001001011101110000010111001100001011010010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33200

pattern = 166; // 33200
ALLPIS = 207'b001100101110010111001110111110110010100011001111101011111110010100001011001101100111010001111000110101110000010000110100100011101000110010000000111000000010000000011010111011010010010101110100110011110110001;
XPCT = 108'b001111010001001010111010011011110110101011111010101110000110000110000101111000010000100110011110010000010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33400

pattern = 167; // 33400
ALLPIS = 207'b110000010100001110001000001001000111111011101110110010111010100100011111000110100110000000100111001010001100010011111110000000100100111111010001011111100110010010000010110011000100100000111000111001111100101;
XPCT = 108'b111110010010010000011100011101111100100011111101111111001111001110001111010111011010111110100001011101010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33600

pattern = 168; // 33600
ALLPIS = 207'b000101101111011010110110011111001001000110000100100111110001010000000110110000001100111001001111011011001001101001100000001001110101011100011001000010010010101011101100110111111110011111011100101100000110110;
XPCT = 108'b000110111111001111101110010100000110101101111010101110000110110101011111010001001001100010011110010111010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33800

pattern = 169; // 33800
ALLPIS = 207'b001110100011110100110001001001000001100111011001111101010111010110101110000100100110101001111001001011010110110001000011101101010110000100100011011101010000010001101011110010001010100110100011101011010000100;
XPCT = 108'b001110010101010011010001110111010000010001101010001010011111001101111111001100001000110111111001000110001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34000

pattern = 170; // 34000
ALLPIS = 207'b000010011011110100110101100010101010111100011100101101100100110110001110101100111001001000010010001101101011110011101001011100100111000010111110110111110000101010101101110110010111000000100001001110001010011;
XPCT = 108'b000110110011100000010000100110001010011101111010001010001111001011000101000111111000111110000000000000000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34200

pattern = 171; // 34200
ALLPIS = 207'b000011000101010101011110101000100110010110100101111001001010010101110001001101010100010100011010001011001101010001100101110000011100110111101101000000100111101010111011100110011000101001110001111010111100111;
XPCT = 108'b001100110100010100111000111110111100011011011010000000001001011100001110001100111011110000100000011000010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34400

pattern = 172; // 34400
ALLPIS = 207'b100000011000001000000010100010100010000100010100110000000000100111000011001010010110100001110101111000111111111000101100110110101110010010110110010010000101011001001010001111011111001110111001100011110001000;
XPCT = 108'b111001110111100111011100110011110001101001101100101111011111101100000101010110100111110010000001011011101110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34600

pattern = 173; // 34600
ALLPIS = 207'b011100100111000010000010010101010010010111110111011110111100100110110100000110110110000110111110100100100000111101101111000000100110110111101100100110110001101001000110010001101110111010101100001011001101111;
XPCT = 108'b001010001111011101010110000111001101100011111001111110001111111111011111011110101011111000011000000000000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34800

pattern = 174; // 34800
ALLPIS = 207'b101001111100101111000001000101101111111001110000111100101001100111010101000010101010111010101010110001000101001110010101101111100001110010111111100111110011010101110011110000011110110100100101010011011000101;
XPCT = 108'b111110000111011010010010101011011000111001111101111111101111110000101111111100100101111111100001100110010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35000

pattern = 175; // 35000
ALLPIS = 207'b100111101000011101010010001111010011100010101011111000100101101100010110110111011010111011000010011011111011001110010010011001001110110111100110011001001011110011100101001110101001111000101101110111011001000;
XPCT = 108'b110001111100111100010110111011011001010101111101011011111001010100001110100100000110110110100001101111101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35200

pattern = 176; // 35200
ALLPIS = 207'b001001001100011111101100000001111100001111000110101010001000110111010111100101100101001010111111110001111011111110000100111001111110101110101000000100001000101101100011010111000111010000101101101100100001000;
XPCT = 108'b001010110011101000010110110100100001110111111001111110011111111110111111100101100110110011100001111011101110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35400

pattern = 177; // 35400
ALLPIS = 207'b000111000000001001100000010100110101010100001110001101011011011101011100110001001111100110111110101100110011101111000100111001111011011011001100111101010110100111111101110101000001110100010111101001000111001;
XPCT = 108'b000110100000111010001011110101000111010000111010001010011001110000101110100101100100111001100001011010100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35600

pattern = 178; // 35600
ALLPIS = 207'b101101100111110100011011010100110101110100100001011010111011101001000100111001000010000000110111011000101100010101111110110100010101101000111011001010101100010001101011000000111011101100111010110001111110000;
XPCT = 108'b111000001101110110011101011001111110111011111100101111011111100100111101000101011111110010011001100010000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35800

pattern = 179; // 35800
ALLPIS = 207'b111110110011000111111000011111000000101110100111011101111111001110000101000101110101110001101010000010111001010010110100010100011001110000110110000010010011010011000000111000100001011101011011011001101100011;
XPCT = 108'b110111001000101110101101101101101100000011111111011011001001111100101110011110110000110001011000001101011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36000

pattern = 180; // 36000
ALLPIS = 207'b011000110010011111001011100001010010011001001000011001000000011000111100001001011111110011111010001110111010010100001001110000001000010001010010111001110010110010010111110100000110110011111011111011010111101;
XPCT = 108'b001110100011011001111101111111010111110011111011111110011111111000001111101101101000111100000000100111100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36200

pattern = 181; // 36200
ALLPIS = 207'b000101010101011101001111100111000111001100110111111000101101010011100111100010111111011111011001011000010000110101001011101111010010100110011001000111000110101111001000000000100101111010101100010011010010101;
XPCT = 108'b000000001010111101010110001011010010100011110000101110001111001000101101111101001001110100111111100111100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36400

pattern = 182; // 36400
ALLPIS = 207'b001101011100100111101110110111011001100100100101011000010000000110010010111101011100001110011010100111011101000111111101110101001100000100111001100101011011010110101000000010010011000010100011011001010000001;
XPCT = 108'b000000010001100001010001101101010000101011111000101110010000010000101010011010001111101111111111011010100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36600

pattern = 183; // 36600
ALLPIS = 207'b011011000101001111010010111111100011100001010010101110100000011111100010000010000001010011101111110010010111011101101011111001001000010001010000110110110110011010011001111000001101001101100011110001001101011;
XPCT = 108'b000111000110100110110001111001001101010011110001011010011001100010101100100101010111111011111000011100011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36800

pattern = 184; // 36800
ALLPIS = 207'b001111000010001111111110010100111000000101001010001001110001101000001000101110010111110000001110001001000111101111011101100101010111111010111101001001000100000111111111110101100001110001111001011110111011100;
XPCT = 108'b001110101000111000111100101110111011010111011010001010000000000001101110001011111000101100111111011011010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37000

pattern = 185; // 37000
ALLPIS = 207'b010001001100011001110100110011001111101100001010111000011001000110110100110111111010001000010110110000100101110011111101001110111001100010100111010110011001110111010110000111111011111010010001110010111111000;
XPCT = 108'b001000111101111101001000111010111111101010111001111110011111010010011111010111001010110111100001000110100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37200

pattern = 186; // 37200
ALLPIS = 207'b110010010111101100001100110000000011100010101000110110000000101000000111100100000111001111100010011000000000110111101011110001001001010110110011100101001110001100000001000010000111011000101110111100100111010;
XPCT = 108'b110000010011101100010111011100100111010111111101011011101111110110101111001111011111111000000111001100110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37400

pattern = 187; // 37400
ALLPIS = 207'b111001110110011111001101100010101100010010000000010001001100101011011011000010010001111110010110001010000110011110011100110000011011100111101101100010001001111110100101000101000001010010101001001000011110101;
XPCT = 108'b110000100000101001010100100100011110110011111111111111101111100101011111101110001100110110100001010111011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37600

pattern = 188; // 37600
ALLPIS = 207'b001111011111011110100001010101100010111011110001111111100010101000010001000010011000001000101111010011100011000111101110111110111110100100001011011111101110101001000100010101010000100110011101010001110111100;
XPCT = 108'b000010100000010011001110101001110111001001111011011010001111101111111111011111111001110110011000001111111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37800

pattern = 189; // 37800
ALLPIS = 207'b000101010101000110101000100110111001100101000111100000011001011010011001001100111010001101001111100011110101111111001110001000010011100011100000111101011010011110011011101100000101010100110110111101101101110;
XPCT = 108'b001101100010101010011011011101101101110111111000101110001001001111001110011100000100111001011000110100010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38000

pattern = 190; // 38000
ALLPIS = 207'b000100001000001001001111000010111101011011001000111011000000010010110101000111100010100111110011101000000111000011100111000110110101100010001110100001110110010110101101010001010111010001100110101100101111000;
XPCT = 108'b000010000011101000110011010100101111111111111010100100001001111111001110000111001001111100100000110000111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38200

pattern = 191; // 38200
ALLPIS = 207'b001101110111101110110110111110001000001100011000101000000110110011000001100110000101110110010100101110001011101001100000010111000001100111000010110101010111111111110000100011111001110110101011110100000110010;
XPCT = 108'b000100011100111011010101111000000110101101111001111110011111100100000101110110111110110100100000100010101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38400

pattern = 192; // 38400
ALLPIS = 207'b100111001000001000000111101001111010000001100101110110110001100110011100001011101111000101101100001011100101110000010000111011110011001100000000010110011101011100001001111000000011010010111011101010011111100;
XPCT = 108'b110111000001101001011101110110011111010001111100001011000110010111101111010000110010101100111111100000111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38600

pattern = 193; // 38600
ALLPIS = 207'b110111100101111110010101110100110001010111110100001001011000011111111010110010000010110000001101010001000101101110100101010100001111111001100101111110000110010101100101101101000011101000010110010110100101000;
XPCT = 108'b110101100001110100001011001010100101010111111111011011011111101011111111100101011011110010011001000110111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38800

pattern = 194; // 38800
ALLPIS = 207'b111001100110001000001000010111001010011101010000001001000000101110001101100001100001000100111010101001110111011000101110010001010100000010101000110000110100100111110111110001100110010101000010001001111100000;
XPCT = 108'b111110001011001010100001000101111100110011111111111111011111011000011111100110100010111011100000010111110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39000

pattern = 195; // 39000
ALLPIS = 207'b110001011000101100010111010110001001001011110111010011010000000100110111110000110110011011101011011110001111010001101010001010101110101110000100000110000101011011010101010010010110000011000110101001010110010;
XPCT = 108'b110010010011000001100011010101010110111011111111111111110000001000001110000011110010100010011001100100101110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39200

pattern = 196; // 39200
ALLPIS = 207'b101101011000001101000000000000110111001011000101011100001001011100010010101011101011010011101101110001110100101101110100100101110111001010100101111010010000001111001010000110000010100001011011000000000110001;
XPCT = 108'b111000110001010000101101100000000110100001111100101111010000100011011110111011111111101110111111001000110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39400

pattern = 197; // 39400
ALLPIS = 207'b001111000000001011010000111010101011010000001001111100101100111111101110100110000010011000110000101110101001000100010111011100010011111101111000110010100001000010011001011011010110010010000100011011101000100;
XPCT = 108'b000011010011001001000010001111101000011001111000001010000000101010111110101010110011101101011111011000101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39600

pattern = 198; // 39600
ALLPIS = 207'b011100010000010111111000011110000101000100001111100101111100101001001001111011101011111100010101100011101101010010001111001011000001000110110010101011110001101101110000011100111100001001000100111001000011101;
XPCT = 108'b000011101110000100100010011101000011101010111011111110010000100111001110110000100001101100111110001100011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39800

pattern = 199; // 39800
ALLPIS = 207'b111011000000111011000111000000101111010011111001000001100001100001101110111010100001000010000010100110001001010110111001001000000010111011110111100000100011001110110110010110011000101100011010010000000111010;
XPCT = 108'b111010110100010110001101001000000111001011111111011011010000011100111100000000001001101101000110000000000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40000

pattern = 200; // 40000
ALLPIS = 207'b010011010001000000011111000111001101100001000101111110100000001000000000110111100100101010011010000000110010000010100100100001101001000011010100001011000111000010111000110011000101000110110111000000100101001;
XPCT = 108'b000110010010100011011011100000100101000011111001011010011111011010001111100110011000110101011110111011000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40200

pattern = 201; // 40200
ALLPIS = 207'b101110010101111101010110010110110001011001100101100000110111011101001111111101111001001101011011100110010100110010010110001101001011010100100110101101001001000101110100100010000010111001011001010010001011001;
XPCT = 108'b110100010001011100101100101010001011000001111101011011111111101110100001010100111110111001011001011100110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40400

pattern = 202; // 40400
ALLPIS = 207'b001101100110000101001000100100001110011111110101111100011000110001110001101101001111100110010110001001101000110000010000100011110111101001100001111111111010111010110011110111011100101001110100101000001000011;
XPCT = 108'b001110110110010100111010010100001000111011111001110100010000111001101110001001001010101011000001111011011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40600

pattern = 203; // 40600
ALLPIS = 207'b110101100011101110111111010111110000101000011110000111101011000001111101111110000110011001100010101000011000111011011001110000101110111101001110000011110110101101011111001010011001111110101001011111000001100;
XPCT = 108'b111001010100111111010100101111000001111111011111111111101111100000001011011111011001111000011000000000011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40800

pattern = 204; // 40800
ALLPIS = 207'b001011011100000001001110101110100101101101011100011000000111101101001110000001010010111111001011011001011110010000001110010001001100011100101000001100111110010111001101101101101010011000011011010000110100110;
XPCT = 108'b000101101101001100001101101000110100010011111000001010000110000111101111100011001000101110011000000111011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41000

pattern = 205; // 41000
ALLPIS = 207'b101100100100010111100011111111011110000110010111001100111111110100001010111011100100010010100110011001001010111101001101111100100000100111101110010100100001111110001110011001010100100110101000000111110100111;
XPCT = 108'b111011000010010011010100000011110100101101111100101111000000111110111110011000100011100111011110010101110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41200

pattern = 206; // 41200
ALLPIS = 207'b101001110000111101101100011110010111010000111001110100100110111110100111110010110001110100000101110001111001000110111110110111010111010101001000110110101000101000110000011011111100101010011100111001111101101;
XPCT = 108'b110011011110010101001110011101111101101011111101111111000000101001011110001011011000100101011111000011100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41400

pattern = 207; // 41400
ALLPIS = 207'b001001011000111100101100011111100101110110101110011100101100010000000001001111001100011101011000111100000001011001011011001111100111111001110010100100010000010001000101110110010000011011111001110111011010011;
XPCT = 108'b000110110000001101111100111011011010111111111001111110010000100100101110001011000010100110000111000010011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41600

pattern = 208; // 41600
ALLPIS = 207'b110011001011011111000101101000110001000001111110111110001001101100110100111000110000011010100100101100011000000011110010111000101010101100101001111111010101000101011010001011111110011100001110001001001111010;
XPCT = 108'b111001011111001110000111000101001111001011111101011011111111100000101111100110001010110100100001101100001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41800

pattern = 209; // 41800
ALLPIS = 207'b100100110011010100000101010000011001010110000101110111010101110110111001101100111111100110100011001001101000111110100101110100000100010100111100011001111001100010010101011001010101101101110110011010100110001;
XPCT = 108'b110011000010110110111011001110100110111001111111110101001111001001011111100100110001110010111111101111010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 42000

pattern = 210; // 42000
ALLPIS = 207'b010011100000001101101100001101011000101111011011010101001011010001111000011110110000011100011000101000101110000110111000011100000110101000100000011011110101010000001101100100010100010101111100110110001001000;
XPCT = 108'b000100100010001010111110011010001001011111111011011010010000000010001110101011011111100000011111001100011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 42200

pattern = 211; // 42200
ALLPIS = 207'b101111011110100101000111000001101001100110001011001101100000110101010111011100010110010101001001000010111011101111001000010000110001000100010111010100110000010001100000101001111001010001101010001100010011111;
XPCT = 108'b110101001100101000110101000100010011001101111111011011000000110011110110011011010100101101011111011000011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 42400

pattern = 212; // 42400
ALLPIS = 207'b011101110010001101111010101110111110111110011110011110010100101110000110000110010011000000111101000111111100010110000110010011001100111100000111111110111100001111101100000110110110000011110100110110011111000;
XPCT = 108'b000000111011000001111010011010011111101111011001111110010110001101001111110011001111101111011110100000000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 42600

pattern = 213; // 42600
ALLPIS = 207'b011000110011101100000111110010111101111111010000100100000001010010011110011110101011000010011000000001101000011100000010101010001001010010011101001100110000000111101010101000110010011010111000000101101111111;
XPCT = 108'b001101001001001101011100000001101111101111111001111110011111111110011111011110000110111001011110010011000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 42800

pattern = 214; // 42800
ALLPIS = 207'b000111010110100100010101011001001001000111101001001010100000001110001111111010000110011110101111100000100010011101001100111000000111000101011111101001100100000111001101110111110100000101101101000110011110011;
XPCT = 108'b000110111010000010110110100010011110011101110000001010010000100111011110010001001111100000100001111011000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 43000

pattern = 215; // 43000
ALLPIS = 207'b100010101000000110000101011010010011011110101110110101011011010110110100001110111001010101010110000111011010100001111100100001110100110011101110101111111010000111110011010110011010100100001001101010110010000;
XPCT = 108'b111010110101010010000100110110110010011001111111010001011111000010001111000100111001110110100000101111111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 43200

pattern = 216; // 43200
ALLPIS = 207'b111110010101000111000010101111001001010110010111010000111111100010001110011101001101101000100100000101110000001101001010011110011100001000100001001110100000011110101011101100110000111101000010110100111111110;
XPCT = 108'b111101101000011110100001011000111111011111111101011011111111000101011111001101000110110001000110101111010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 43400

pattern = 217; // 43400
ALLPIS = 207'b100100000111111111101000011000110000000010100011011111101100110000011110110111101111011100010111110100000100101010001000001010001001010011100000001101111000000000000001111001001111110001001100010101000100001;
XPCT = 108'b110111000111111000100110001001000100110111111111111111111111101111111111100111100000111011111111000010101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 43600

pattern = 218; // 43600
ALLPIS = 207'b110000011100101011011010101101011000001001110110101001001100011100110101100000000101011000101111111011010110111011100011110010111001111010111100101000110110110001111100110010101001010000110101000111101101110;
XPCT = 108'b110110011100101000011010100011101101100111101111111111110000100000011110010000101000101101011000110111110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 43800

pattern = 219; // 43800
ALLPIS = 207'b010110010001111100100011011000110010111011110101000111000111100011101000101111111010111011100110110100010101010111101100011000010110111110111100110001011011101000010001100001001100111010000110001100111110000;
XPCT = 108'b000100000110011101000011000100111110010111111011011010001111001010100101000110011100111000111111011110001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 44000

pattern = 220; // 44000
ALLPIS = 207'b010100011010100110000111011010010100100100011011001111001110101110111000001010011111100011010010011111100001011010110110100100101011001011100101101000001100000111101010110101111010000101111010110010100101101;
XPCT = 108'b001110101101000010111101011010100101101011111011111110001111010000011111010101101000110111000000000101101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 44200

pattern = 221; // 44200
ALLPIS = 207'b000111110111101101111110101010011001001101010010110101011010011101110000011001100000111010110111011000010101000011100111111010001010100100100111001001100111111110001001010010100100011000110011100101100100110;
XPCT = 108'b000010011010001100011001110001100100010111111010000000001001101110001110111111101011111111100000010101011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 44400

pattern = 222; // 44400
ALLPIS = 207'b100101011110011000101110000100011100000011110011011111010110101001111011011010100110100000111110101000101011000011100010100110100010011101000001110100010110110110011110001011001000010011000010111001000111001;
XPCT = 108'b111001010100001001100001011101000111100010111110100101010000010111101110001001011010101000111110001100101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 44600

pattern = 223; // 44600
ALLPIS = 207'b000100100110001000100100111010000100000001101000011110100110111011110100100111000110100100011000110010010010010001000011011111001100101011101110111100001101011011000111001111100000111110101001010001010011110;
XPCT = 108'b001001111000011111010100101001010011110001111001110100000110011100011111000010010111100000100110101011111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 44800

pattern = 224; // 44800
ALLPIS = 207'b000000100001001000111101110110000111001011000111111011000100010011010010000100100111011010111000001001110110101001001111001010011011100110100101101110100001111000011101011100110110011011100001000110000101100;
XPCT = 108'b000011101011001101110000100010000101111111111010101110011111101000011111001100010001111001011111010011000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 45000

pattern = 225; // 45000
ALLPIS = 207'b011000111010101110101101010010110101010010100110010110000010010010101000011100010110110111111000110001010000101010010110110011111101101111000100111110010100101010000001110100001000001001100111001110011010111;
XPCT = 108'b000110100100000100110011100110011010110111111001111110000000011001111110001010111010101011011110001000011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 45200

pattern = 226; // 45200
ALLPIS = 207'b000101100111110011101100001001111000010101010101010100011011110010000001001100001111010111111110001011001111001111111000101000001111101111110100100011100101100000100000001101010110010001011000000100011111110;
XPCT = 108'b000001100011001000101100000000011111101111111001111110001111101001011111101110000111111110111001010001001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 45400

pattern = 227; // 45400
ALLPIS = 207'b110101100001001110110000101011011110101010010011100001110001111010000010111101011000110000011001000111001101111100110001101110100111111110111000001101110110110110101011100000100011100011101000111111001100011;
XPCT = 108'b111100001001110001110100011111001100110111110111111111011001000011111110000111001000110011111111001110110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 45600

pattern = 228; // 45600
ALLPIS = 207'b111001110000111101010001100010111110101110100010011110000000011110101011001110111011001100001101111001100000010100111010011011000110011011111101010110101000010001010010011010100010001100100001101001011100111;
XPCT = 108'b111011011001000110010000110101011100100011111101111111100000000010111110111001110010101111011001100000110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 45800

pattern = 229; // 45800
ALLPIS = 207'b101000100000111011000001110000111001101010001011111101111000000100010100001000000101000001101101010011011001110001011000100001100111011100011111010111101011100110110111001100000110110010111101100101010111110;
XPCT = 108'b111001100011011001011110110001010111110101111111111111010000010101011110100000100101101100111110000001011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 46000

pattern = 230; // 46000
ALLPIS = 207'b010110111000010110010101100001111101110001111000001110000000100001000000110010011010011000111010000001111000011011110001111001100101110000011110100110010110011001110110100010100010101100001000101110110101001;
XPCT = 108'b001100011001010110000100010110110101000111111001011010011111101001011111111101001110110010100000011000101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 46200

pattern = 231; // 46200
ALLPIS = 207'b011110011011111001101011101111111010000001110100101101101111111001110100111110010010110110111010101001111000110010010101111000001100001110101101001000111110101011011000110000000010101111001001000111101110101;
XPCT = 108'b000110000001010111100100100011101110000111111011011010001111111101101111111111011000110010011000110001000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 46400

pattern = 232; // 46400
ALLPIS = 207'b000010001011101001111001100101000011100000000110111011100010001001011000011010010101000101001010010001111001011010110100100000010011011100001001110100001111010100001000100101101011100111110011011000111000000;
XPCT = 108'b000100101101110011111001101100111000000011111010001010011111010101101011011111111100110101111110010100010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 46600

pattern = 233; // 46600
ALLPIS = 207'b101111010001010000011011000111100010011101100010100111000010111000011000110010011111001100110010111100000111001011001111110110111001010111010110000100011001111001011111111111011000100101011110110111110011011;
XPCT = 108'b111111110100010010101111011011110011011110111110001011110110101010011111000001010000100111011110100101101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 46800

pattern = 234; // 46800
ALLPIS = 207'b111000011000001100010011000101100010101010010001001010000000000111111000111110001111100000110110011101011101100000010101001000101101100111000101001001111000101000100101100011000101110010100011000110100010100;
XPCT = 108'b110100010010111001010001100010100010110111111101111111001111101001001111100100101110111100100000011100010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 47000

pattern = 235; // 47000
ALLPIS = 207'b110000101110011001111010111010101100100010000111001000100111000001110111111100110111111001110110111100101111001011011010111011001111000001101010010100101001011000010001100100101010111011001001011111101001110;
XPCT = 108'b110100101101011101100100101111101001110111111101111111110000000001111110000001101110101000011110001101000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 47200

pattern = 236; // 47200
ALLPIS = 207'b100010100101110001000100100011100101001100010000011110111011011101011101011001010001110110011111100000001000101010101110001111010000100001101001001001011110100000100111100100110011001000111101001100001101101;
XPCT = 108'b111100101001100100011110100100001101011101111101011011011111110110101111000100101110111011011110111111110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 47400

pattern = 237; // 47400
ALLPIS = 207'b011110100011100100010011011011000000111011001100000111001010000100011111111101011100111100010001101110000111111111000011001000000011000111001100111101010001110000110111100000100111100101111111111100011111011;
XPCT = 108'b001100001011110010111111111100011111010110100011011010011111110011000001001110011100110110011000111110110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 47600

pattern = 238; // 47600
ALLPIS = 207'b010000110010111000110100001110011001011000011010111011110110100101000110011110101011000111011111001001101111111011001101010110110010010011000101010100110111000100110101001011110010101011100110100111110110111;
XPCT = 108'b000001011001010101110011010011110110111110001011111110000110010100000001000001000101101010111001011101000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 47800

pattern = 239; // 47800
ALLPIS = 207'b010010100100111111001110110111101111100111000000111101111000111010101011111100010110111111100111100101010111010101000011111100000100111100110101110011010100101111111011001110010101011111100110011010110100111;
XPCT = 108'b001001110010101111110011001110110100011010010011011010000000101100000000001001000101100001100110010110010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 48000

pattern = 240; // 48000
ALLPIS = 207'b001100011110011010101000101111100010000000111001111111011110111010001100111000010011101011111000100001000111010111010110011000110001001000101111100011110011110011101011110011101110101001011100110111011001001;
XPCT = 108'b001110011111010100101110011011011001110111111010101110000000110011011110100011101000101010111110011001010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 48200

      $display("// %t : Simulation of %0d patterns completed with %0d errors\n", $time, pattern+1, nofails);
      if (verbose >=2) $finish(2);
      /* else */ $finish(0);
   end
endmodule
