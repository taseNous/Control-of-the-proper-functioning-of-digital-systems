// Verilog pattern output written by  TetraMAX (TM)  B-2008.09-SP2-i081128_181834 
// Date: Wed Jul  6 12:08:39 2011
// Module tested: c7552

//     Uncollapsed Stuck Fault Summary Report
// -----------------------------------------------
// fault class                     code   #faults
// ------------------------------  ----  ---------
// Detected                         DT       6122
// Possibly detected                PT          0
// Undetectable                     UD          0
// ATPG untestable                  AU          0
// Not detected                     ND        766
// -----------------------------------------------
// total faults                              6888
// test coverage                            88.88%
// -----------------------------------------------
// 
//            Pattern Summary Report
// -----------------------------------------------
// #internal patterns                          77
//     #basic_scan patterns                    77
// -----------------------------------------------
// 
// There are no rule fails
// There are no clocks
// There are no constraint ports
// There are no equivalent pins
// There are no net connections

`timescale 1 ns / 1 ns

//
// --- NOTE: Remove the comment to define 'tmax_iddq' to activate processing of IDDQ events
//     Or use '+define+tmax_iddq' on the verilog compile line
//
//`define tmax_iddq

module AAA_tmax_testbench_1_16 ;
   parameter NAMELENGTH = 200; // max length of names reported in fails
   integer nofails, bit, pattern, lastpattern;
   integer error_banner; // flag for tracking displayed error banner
   integer loads;        // number of load_unloads for current pattern
   integer patm1;        // pattern - 1
   integer patp1;        // pattern + lastpattern
   integer prev_pat;     // previous pattern number
   integer report_interval; // report pattern progress every Nth pattern
   integer verbose;      // message verbosity level
   parameter NINPUTS = 207, NOUTPUTS = 108;
   wire [0:NOUTPUTS-1] PO; reg [0:NOUTPUTS-1] ALLPOS, XPCT, MASK;
   reg [0:NINPUTS-1] PI, ALLPIS;
   reg [0:8*(NAMELENGTH-1)] POnames [0:NOUTPUTS-1];
   event IDDQ;

   wire N1;
   wire N5;
   wire N9;
   wire N12;
   wire N15;
   wire N18;
   wire N23;
   wire N26;
   wire N29;
   wire N32;
   wire N35;
   wire N38;
   wire N41;
   wire N44;
   wire N47;
   wire N50;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N69;
   wire N70;
   wire N73;
   wire N74;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N82;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N94;
   wire N97;
   wire N100;
   wire N103;
   wire N106;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N118;
   wire N121;
   wire N124;
   wire N127;
   wire N130;
   wire N133;
   wire N134;
   wire N135;
   wire N138;
   wire N141;
   wire N144;
   wire N147;
   wire N150;
   wire N151;
   wire N152;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N178;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire N185;
   wire N186;
   wire N187;
   wire N188;
   wire N189;
   wire N190;
   wire N191;
   wire N192;
   wire N193;
   wire N194;
   wire N195;
   wire N196;
   wire N197;
   wire N198;
   wire N199;
   wire N200;
   wire N201;
   wire N202;
   wire N203;
   wire N204;
   wire N205;
   wire N206;
   wire N207;
   wire N208;
   wire N209;
   wire N210;
   wire N211;
   wire N212;
   wire N213;
   wire N214;
   wire N215;
   wire N216;
   wire N217;
   wire N218;
   wire N219;
   wire N220;
   wire N221;
   wire N222;
   wire N223;
   wire N224;
   wire N225;
   wire N226;
   wire N227;
   wire N228;
   wire N229;
   wire N230;
   wire N231;
   wire N232;
   wire N233;
   wire N234;
   wire N235;
   wire N236;
   wire N237;
   wire N238;
   wire N239;
   wire N240;
   wire N242;
   wire N245;
   wire N248;
   wire N251;
   wire N254;
   wire N257;
   wire N260;
   wire N263;
   wire N267;
   wire N271;
   wire N274;
   wire N277;
   wire N280;
   wire N283;
   wire N286;
   wire N289;
   wire N293;
   wire N296;
   wire N299;
   wire N303;
   wire N307;
   wire N310;
   wire N313;
   wire N316;
   wire N319;
   wire N322;
   wire N325;
   wire N328;
   wire N331;
   wire N334;
   wire N337;
   wire N340;
   wire N343;
   wire N346;
   wire N349;
   wire N352;
   wire N355;
   wire N358;
   wire N361;
   wire N364;
   wire N367;
   wire N382;
   wire N241_I;
   wire N387;
   wire N388;
   wire N478;
   wire N482;
   wire N484;
   wire N486;
   wire N489;
   wire N492;
   wire N501;
   wire N505;
   wire N507;
   wire N509;
   wire N511;
   wire N513;
   wire N515;
   wire N517;
   wire N519;
   wire N535;
   wire N537;
   wire N539;
   wire N541;
   wire N543;
   wire N545;
   wire N547;
   wire N549;
   wire N551;
   wire N553;
   wire N556;
   wire N559;
   wire N561;
   wire N563;
   wire N565;
   wire N567;
   wire N569;
   wire N571;
   wire N573;
   wire N582;
   wire N643;
   wire N707;
   wire N813;
   wire N881;
   wire N882;
   wire N883;
   wire N884;
   wire N885;
   wire N889;
   wire N945;
   wire N1110;
   wire N1111;
   wire N1112;
   wire N1113;
   wire N1114;
   wire N1489;
   wire N1490;
   wire N1781;
   wire N10025;
   wire N10101;
   wire N10102;
   wire N10103;
   wire N10104;
   wire N10109;
   wire N10110;
   wire N10111;
   wire N10112;
   wire N10350;
   wire N10351;
   wire N10352;
   wire N10353;
   wire N10574;
   wire N10575;
   wire N10576;
   wire N10628;
   wire N10632;
   wire N10641;
   wire N10704;
   wire N10706;
   wire N10711;
   wire N10712;
   wire N10713;
   wire N10714;
   wire N10715;
   wire N10716;
   wire N10717;
   wire N10718;
   wire N10729;
   wire N10759;
   wire N10760;
   wire N10761;
   wire N10762;
   wire N10763;
   wire N10827;
   wire N10837;
   wire N10838;
   wire N10839;
   wire N10840;
   wire N10868;
   wire N10869;
   wire N10870;
   wire N10871;
   wire N10905;
   wire N10906;
   wire N10907;
   wire N10908;
   wire N11333;
   wire N11334;
   wire N11340;
   wire N11342;
   wire N241_O;

   // map PI[] vector to DUT inputs and bidis
   assign N1 = PI[0];
   assign N5 = PI[1];
   assign N9 = PI[2];
   assign N12 = PI[3];
   assign N15 = PI[4];
   assign N18 = PI[5];
   assign N23 = PI[6];
   assign N26 = PI[7];
   assign N29 = PI[8];
   assign N32 = PI[9];
   assign N35 = PI[10];
   assign N38 = PI[11];
   assign N41 = PI[12];
   assign N44 = PI[13];
   assign N47 = PI[14];
   assign N50 = PI[15];
   assign N53 = PI[16];
   assign N54 = PI[17];
   assign N55 = PI[18];
   assign N56 = PI[19];
   assign N57 = PI[20];
   assign N58 = PI[21];
   assign N59 = PI[22];
   assign N60 = PI[23];
   assign N61 = PI[24];
   assign N62 = PI[25];
   assign N63 = PI[26];
   assign N64 = PI[27];
   assign N65 = PI[28];
   assign N66 = PI[29];
   assign N69 = PI[30];
   assign N70 = PI[31];
   assign N73 = PI[32];
   assign N74 = PI[33];
   assign N75 = PI[34];
   assign N76 = PI[35];
   assign N77 = PI[36];
   assign N78 = PI[37];
   assign N79 = PI[38];
   assign N80 = PI[39];
   assign N81 = PI[40];
   assign N82 = PI[41];
   assign N83 = PI[42];
   assign N84 = PI[43];
   assign N85 = PI[44];
   assign N86 = PI[45];
   assign N87 = PI[46];
   assign N88 = PI[47];
   assign N89 = PI[48];
   assign N94 = PI[49];
   assign N97 = PI[50];
   assign N100 = PI[51];
   assign N103 = PI[52];
   assign N106 = PI[53];
   assign N109 = PI[54];
   assign N110 = PI[55];
   assign N111 = PI[56];
   assign N112 = PI[57];
   assign N113 = PI[58];
   assign N114 = PI[59];
   assign N115 = PI[60];
   assign N118 = PI[61];
   assign N121 = PI[62];
   assign N124 = PI[63];
   assign N127 = PI[64];
   assign N130 = PI[65];
   assign N133 = PI[66];
   assign N134 = PI[67];
   assign N135 = PI[68];
   assign N138 = PI[69];
   assign N141 = PI[70];
   assign N144 = PI[71];
   assign N147 = PI[72];
   assign N150 = PI[73];
   assign N151 = PI[74];
   assign N152 = PI[75];
   assign N153 = PI[76];
   assign N154 = PI[77];
   assign N155 = PI[78];
   assign N156 = PI[79];
   assign N157 = PI[80];
   assign N158 = PI[81];
   assign N159 = PI[82];
   assign N160 = PI[83];
   assign N161 = PI[84];
   assign N162 = PI[85];
   assign N163 = PI[86];
   assign N164 = PI[87];
   assign N165 = PI[88];
   assign N166 = PI[89];
   assign N167 = PI[90];
   assign N168 = PI[91];
   assign N169 = PI[92];
   assign N170 = PI[93];
   assign N171 = PI[94];
   assign N172 = PI[95];
   assign N173 = PI[96];
   assign N174 = PI[97];
   assign N175 = PI[98];
   assign N176 = PI[99];
   assign N177 = PI[100];
   assign N178 = PI[101];
   assign N179 = PI[102];
   assign N180 = PI[103];
   assign N181 = PI[104];
   assign N182 = PI[105];
   assign N183 = PI[106];
   assign N184 = PI[107];
   assign N185 = PI[108];
   assign N186 = PI[109];
   assign N187 = PI[110];
   assign N188 = PI[111];
   assign N189 = PI[112];
   assign N190 = PI[113];
   assign N191 = PI[114];
   assign N192 = PI[115];
   assign N193 = PI[116];
   assign N194 = PI[117];
   assign N195 = PI[118];
   assign N196 = PI[119];
   assign N197 = PI[120];
   assign N198 = PI[121];
   assign N199 = PI[122];
   assign N200 = PI[123];
   assign N201 = PI[124];
   assign N202 = PI[125];
   assign N203 = PI[126];
   assign N204 = PI[127];
   assign N205 = PI[128];
   assign N206 = PI[129];
   assign N207 = PI[130];
   assign N208 = PI[131];
   assign N209 = PI[132];
   assign N210 = PI[133];
   assign N211 = PI[134];
   assign N212 = PI[135];
   assign N213 = PI[136];
   assign N214 = PI[137];
   assign N215 = PI[138];
   assign N216 = PI[139];
   assign N217 = PI[140];
   assign N218 = PI[141];
   assign N219 = PI[142];
   assign N220 = PI[143];
   assign N221 = PI[144];
   assign N222 = PI[145];
   assign N223 = PI[146];
   assign N224 = PI[147];
   assign N225 = PI[148];
   assign N226 = PI[149];
   assign N227 = PI[150];
   assign N228 = PI[151];
   assign N229 = PI[152];
   assign N230 = PI[153];
   assign N231 = PI[154];
   assign N232 = PI[155];
   assign N233 = PI[156];
   assign N234 = PI[157];
   assign N235 = PI[158];
   assign N236 = PI[159];
   assign N237 = PI[160];
   assign N238 = PI[161];
   assign N239 = PI[162];
   assign N240 = PI[163];
   assign N242 = PI[164];
   assign N245 = PI[165];
   assign N248 = PI[166];
   assign N251 = PI[167];
   assign N254 = PI[168];
   assign N257 = PI[169];
   assign N260 = PI[170];
   assign N263 = PI[171];
   assign N267 = PI[172];
   assign N271 = PI[173];
   assign N274 = PI[174];
   assign N277 = PI[175];
   assign N280 = PI[176];
   assign N283 = PI[177];
   assign N286 = PI[178];
   assign N289 = PI[179];
   assign N293 = PI[180];
   assign N296 = PI[181];
   assign N299 = PI[182];
   assign N303 = PI[183];
   assign N307 = PI[184];
   assign N310 = PI[185];
   assign N313 = PI[186];
   assign N316 = PI[187];
   assign N319 = PI[188];
   assign N322 = PI[189];
   assign N325 = PI[190];
   assign N328 = PI[191];
   assign N331 = PI[192];
   assign N334 = PI[193];
   assign N337 = PI[194];
   assign N340 = PI[195];
   assign N343 = PI[196];
   assign N346 = PI[197];
   assign N349 = PI[198];
   assign N352 = PI[199];
   assign N355 = PI[200];
   assign N358 = PI[201];
   assign N361 = PI[202];
   assign N364 = PI[203];
   assign N367 = PI[204];
   assign N382 = PI[205];
   assign N241_I = PI[206];

   // map DUT outputs and bidis to PO[] vector
   assign
      PO[0] = N387 ,
      PO[1] = N388 ,
      PO[2] = N478 ,
      PO[3] = N482 ,
      PO[4] = N484 ,
      PO[5] = N486 ,
      PO[6] = N489 ,
      PO[7] = N492 ,
      PO[8] = N501 ,
      PO[9] = N505 ,
      PO[10] = N507 ,
      PO[11] = N509 ,
      PO[12] = N511 ,
      PO[13] = N513 ,
      PO[14] = N515 ,
      PO[15] = N517 ,
      PO[16] = N519 ,
      PO[17] = N535 ,
      PO[18] = N537 ,
      PO[19] = N539 ,
      PO[20] = N541 ,
      PO[21] = N543 ,
      PO[22] = N545 ,
      PO[23] = N547 ,
      PO[24] = N549 ,
      PO[25] = N551 ,
      PO[26] = N553 ,
      PO[27] = N556 ,
      PO[28] = N559 ,
      PO[29] = N561 ,
      PO[30] = N563 ,
      PO[31] = N565 ;
   assign
      PO[32] = N567 ,
      PO[33] = N569 ,
      PO[34] = N571 ,
      PO[35] = N573 ,
      PO[36] = N582 ,
      PO[37] = N643 ,
      PO[38] = N707 ,
      PO[39] = N813 ,
      PO[40] = N881 ,
      PO[41] = N882 ,
      PO[42] = N883 ,
      PO[43] = N884 ,
      PO[44] = N885 ,
      PO[45] = N889 ,
      PO[46] = N945 ,
      PO[47] = N1110 ,
      PO[48] = N1111 ,
      PO[49] = N1112 ,
      PO[50] = N1113 ,
      PO[51] = N1114 ,
      PO[52] = N1489 ,
      PO[53] = N1490 ,
      PO[54] = N1781 ,
      PO[55] = N10025 ,
      PO[56] = N10101 ,
      PO[57] = N10102 ,
      PO[58] = N10103 ,
      PO[59] = N10104 ,
      PO[60] = N10109 ,
      PO[61] = N10110 ,
      PO[62] = N10111 ,
      PO[63] = N10112 ;
   assign
      PO[64] = N10350 ,
      PO[65] = N10351 ,
      PO[66] = N10352 ,
      PO[67] = N10353 ,
      PO[68] = N10574 ,
      PO[69] = N10575 ,
      PO[70] = N10576 ,
      PO[71] = N10628 ,
      PO[72] = N10632 ,
      PO[73] = N10641 ,
      PO[74] = N10704 ,
      PO[75] = N10706 ,
      PO[76] = N10711 ,
      PO[77] = N10712 ,
      PO[78] = N10713 ,
      PO[79] = N10714 ,
      PO[80] = N10715 ,
      PO[81] = N10716 ,
      PO[82] = N10717 ,
      PO[83] = N10718 ,
      PO[84] = N10729 ,
      PO[85] = N10759 ,
      PO[86] = N10760 ,
      PO[87] = N10761 ,
      PO[88] = N10762 ,
      PO[89] = N10763 ,
      PO[90] = N10827 ,
      PO[91] = N10837 ,
      PO[92] = N10838 ,
      PO[93] = N10839 ,
      PO[94] = N10840 ,
      PO[95] = N10868 ;
   assign
      PO[96] = N10869 ,
      PO[97] = N10870 ,
      PO[98] = N10871 ,
      PO[99] = N10905 ,
      PO[100] = N10906 ,
      PO[101] = N10907 ,
      PO[102] = N10908 ,
      PO[103] = N11333 ,
      PO[104] = N11334 ,
      PO[105] = N11340 ,
      PO[106] = N11342 ,
      PO[107] = N241_O ;

   // instantiate the design into the testbench
   c7552 dut (
      .N1(N1),
      .N5(N5),
      .N9(N9),
      .N12(N12),
      .N15(N15),
      .N18(N18),
      .N23(N23),
      .N26(N26),
      .N29(N29),
      .N32(N32),
      .N35(N35),
      .N38(N38),
      .N41(N41),
      .N44(N44),
      .N47(N47),
      .N50(N50),
      .N53(N53),
      .N54(N54),
      .N55(N55),
      .N56(N56),
      .N57(N57),
      .N58(N58),
      .N59(N59),
      .N60(N60),
      .N61(N61),
      .N62(N62),
      .N63(N63),
      .N64(N64),
      .N65(N65),
      .N66(N66),
      .N69(N69),
      .N70(N70),
      .N73(N73),
      .N74(N74),
      .N75(N75),
      .N76(N76),
      .N77(N77),
      .N78(N78),
      .N79(N79),
      .N80(N80),
      .N81(N81),
      .N82(N82),
      .N83(N83),
      .N84(N84),
      .N85(N85),
      .N86(N86),
      .N87(N87),
      .N88(N88),
      .N89(N89),
      .N94(N94),
      .N97(N97),
      .N100(N100),
      .N103(N103),
      .N106(N106),
      .N109(N109),
      .N110(N110),
      .N111(N111),
      .N112(N112),
      .N113(N113),
      .N114(N114),
      .N115(N115),
      .N118(N118),
      .N121(N121),
      .N124(N124),
      .N127(N127),
      .N130(N130),
      .N133(N133),
      .N134(N134),
      .N135(N135),
      .N138(N138),
      .N141(N141),
      .N144(N144),
      .N147(N147),
      .N150(N150),
      .N151(N151),
      .N152(N152),
      .N153(N153),
      .N154(N154),
      .N155(N155),
      .N156(N156),
      .N157(N157),
      .N158(N158),
      .N159(N159),
      .N160(N160),
      .N161(N161),
      .N162(N162),
      .N163(N163),
      .N164(N164),
      .N165(N165),
      .N166(N166),
      .N167(N167),
      .N168(N168),
      .N169(N169),
      .N170(N170),
      .N171(N171),
      .N172(N172),
      .N173(N173),
      .N174(N174),
      .N175(N175),
      .N176(N176),
      .N177(N177),
      .N178(N178),
      .N179(N179),
      .N180(N180),
      .N181(N181),
      .N182(N182),
      .N183(N183),
      .N184(N184),
      .N185(N185),
      .N186(N186),
      .N187(N187),
      .N188(N188),
      .N189(N189),
      .N190(N190),
      .N191(N191),
      .N192(N192),
      .N193(N193),
      .N194(N194),
      .N195(N195),
      .N196(N196),
      .N197(N197),
      .N198(N198),
      .N199(N199),
      .N200(N200),
      .N201(N201),
      .N202(N202),
      .N203(N203),
      .N204(N204),
      .N205(N205),
      .N206(N206),
      .N207(N207),
      .N208(N208),
      .N209(N209),
      .N210(N210),
      .N211(N211),
      .N212(N212),
      .N213(N213),
      .N214(N214),
      .N215(N215),
      .N216(N216),
      .N217(N217),
      .N218(N218),
      .N219(N219),
      .N220(N220),
      .N221(N221),
      .N222(N222),
      .N223(N223),
      .N224(N224),
      .N225(N225),
      .N226(N226),
      .N227(N227),
      .N228(N228),
      .N229(N229),
      .N230(N230),
      .N231(N231),
      .N232(N232),
      .N233(N233),
      .N234(N234),
      .N235(N235),
      .N236(N236),
      .N237(N237),
      .N238(N238),
      .N239(N239),
      .N240(N240),
      .N242(N242),
      .N245(N245),
      .N248(N248),
      .N251(N251),
      .N254(N254),
      .N257(N257),
      .N260(N260),
      .N263(N263),
      .N267(N267),
      .N271(N271),
      .N274(N274),
      .N277(N277),
      .N280(N280),
      .N283(N283),
      .N286(N286),
      .N289(N289),
      .N293(N293),
      .N296(N296),
      .N299(N299),
      .N303(N303),
      .N307(N307),
      .N310(N310),
      .N313(N313),
      .N316(N316),
      .N319(N319),
      .N322(N322),
      .N325(N325),
      .N328(N328),
      .N331(N331),
      .N334(N334),
      .N337(N337),
      .N340(N340),
      .N343(N343),
      .N346(N346),
      .N349(N349),
      .N352(N352),
      .N355(N355),
      .N358(N358),
      .N361(N361),
      .N364(N364),
      .N367(N367),
      .N382(N382),
      .N241_I(N241_I),
      .N387(N387),
      .N388(N388),
      .N478(N478),
      .N482(N482),
      .N484(N484),
      .N486(N486),
      .N489(N489),
      .N492(N492),
      .N501(N501),
      .N505(N505),
      .N507(N507),
      .N509(N509),
      .N511(N511),
      .N513(N513),
      .N515(N515),
      .N517(N517),
      .N519(N519),
      .N535(N535),
      .N537(N537),
      .N539(N539),
      .N541(N541),
      .N543(N543),
      .N545(N545),
      .N547(N547),
      .N549(N549),
      .N551(N551),
      .N553(N553),
      .N556(N556),
      .N559(N559),
      .N561(N561),
      .N563(N563),
      .N565(N565),
      .N567(N567),
      .N569(N569),
      .N571(N571),
      .N573(N573),
      .N582(N582),
      .N643(N643),
      .N707(N707),
      .N813(N813),
      .N881(N881),
      .N882(N882),
      .N883(N883),
      .N884(N884),
      .N885(N885),
      .N889(N889),
      .N945(N945),
      .N1110(N1110),
      .N1111(N1111),
      .N1112(N1112),
      .N1113(N1113),
      .N1114(N1114),
      .N1489(N1489),
      .N1490(N1490),
      .N1781(N1781),
      .N10025(N10025),
      .N10101(N10101),
      .N10102(N10102),
      .N10103(N10103),
      .N10104(N10104),
      .N10109(N10109),
      .N10110(N10110),
      .N10111(N10111),
      .N10112(N10112),
      .N10350(N10350),
      .N10351(N10351),
      .N10352(N10352),
      .N10353(N10353),
      .N10574(N10574),
      .N10575(N10575),
      .N10576(N10576),
      .N10628(N10628),
      .N10632(N10632),
      .N10641(N10641),
      .N10704(N10704),
      .N10706(N10706),
      .N10711(N10711),
      .N10712(N10712),
      .N10713(N10713),
      .N10714(N10714),
      .N10715(N10715),
      .N10716(N10716),
      .N10717(N10717),
      .N10718(N10718),
      .N10729(N10729),
      .N10759(N10759),
      .N10760(N10760),
      .N10761(N10761),
      .N10762(N10762),
      .N10763(N10763),
      .N10827(N10827),
      .N10837(N10837),
      .N10838(N10838),
      .N10839(N10839),
      .N10840(N10840),
      .N10868(N10868),
      .N10869(N10869),
      .N10870(N10870),
      .N10871(N10871),
      .N10905(N10905),
      .N10906(N10906),
      .N10907(N10907),
      .N10908(N10908),
      .N11333(N11333),
      .N11334(N11334),
      .N11340(N11340),
      .N11342(N11342),
      .N241_O(N241_O)   );


   integer errshown;
   event measurePO;
   always @ measurePO begin
      if (((XPCT&MASK) !== (ALLPOS&MASK)) || (XPCT !== (~(~XPCT)))) begin
         errshown = 0;
         for (bit = 0; bit < NOUTPUTS; bit=bit + 1) begin
            if (MASK[bit]==1'b1) begin
               if (XPCT[bit] !== ALLPOS[bit]) begin
                  if (errshown==0) $display("\n// *** ERROR during capture pattern %0d, T=%t", pattern, $time);
                  $display("  %0d %0s (exp=%b, got=%b)", pattern, POnames[bit], XPCT[bit], ALLPOS[bit]);
                  nofails = nofails + 1; errshown = 1;
               end
            end
         end
      end
   end

   event forcePI_default_WFT;
   always @ forcePI_default_WFT begin
      PI = ALLPIS;
   end
   event measurePO_default_WFT;
   always @ measurePO_default_WFT begin
      #40;
      ALLPOS = PO;
      #0; #0 -> measurePO;
      `ifdef tmax_iddq
         #0; ->IDDQ;
      `endif
   end

   always @ IDDQ begin
   `ifdef tmax_iddq
      $ssi_iddq("strobe_try");
      $ssi_iddq("status drivers leaky AAA_tmax_testbench_1_16.leaky");
   `endif
   end

   event capture;
   always @ capture begin
      ->forcePI_default_WFT;
      #100; ->measurePO_default_WFT;
   end


   initial begin

      //
      // --- establish a default time format for %t
      //
      $timeformat(-9,2," ns",18);

      //
      // --- default verbosity to 2 but also allow user override by
      //     using '+define+tmax_msg=N' on verilog compile line.
      //
      `ifdef tmax_msg
         verbose = `tmax_msg ;
      `else
         verbose = 2 ;
      `endif

      //
      // --- default pattern reporting interval to 5 but also allow user
      //     override by using '+define+tmax_rpt=N' on verilog compile line.
      //
      `ifdef tmax_rpt
         report_interval = `tmax_rpt ;
      `else
         report_interval = 5 ;
      `endif

      //
      // --- support generating Extened VCD output by using
      //     '+define+tmax_vcde' on verilog compile line.
      //
      `ifdef tmax_vcde
         // extended VCD, see IEEE Verilog P1364.1-1999 Draft 2
         if (verbose >= 2) $display("// %t : opening Extended VCD output file", $time);
         $dumpports( dut, "sim_vcde.out");
      `endif

      //
      // --- IDDQ PLI initialization
      //     User may activite by using '+define+tmax_iddq' on verilog compile line.
      //     Or by defining `tmax_iddq in this file.
      //
      `ifdef tmax_iddq
         if (verbose >= 3) $display("// %t : Initializing IDDQ PLI", $time);
         $ssi_iddq("dut AAA_tmax_testbench_1_16.dut");
         $ssi_iddq("verb on");
         $ssi_iddq("cycle 0");
         //
         // --- User may select one of the following two methods for fault seeding:
         //     #1 faults seeded by PLI (default)
         //     #2 faults supplied in a file
         //     Comment out the unused lines as needed (precede with '//').
         //     Replace the 'FAULTLIST_FILE' string with the actual file pathname.
         //
         $ssi_iddq("seed SA AAA_tmax_testbench_1_16.dut");   // no file, faults seeded by PLI
         //
         // $ssi_iddq("scope AAA_tmax_testbench_1_16.dut");   // set scope for faults from a file
         // $ssi_iddq("read_tmax FAULTLIST_FILE"); // read faults from a file
         //
      `endif

      POnames[0] = "N387";
      POnames[1] = "N388";
      POnames[2] = "N478";
      POnames[3] = "N482";
      POnames[4] = "N484";
      POnames[5] = "N486";
      POnames[6] = "N489";
      POnames[7] = "N492";
      POnames[8] = "N501";
      POnames[9] = "N505";
      POnames[10] = "N507";
      POnames[11] = "N509";
      POnames[12] = "N511";
      POnames[13] = "N513";
      POnames[14] = "N515";
      POnames[15] = "N517";
      POnames[16] = "N519";
      POnames[17] = "N535";
      POnames[18] = "N537";
      POnames[19] = "N539";
      POnames[20] = "N541";
      POnames[21] = "N543";
      POnames[22] = "N545";
      POnames[23] = "N547";
      POnames[24] = "N549";
      POnames[25] = "N551";
      POnames[26] = "N553";
      POnames[27] = "N556";
      POnames[28] = "N559";
      POnames[29] = "N561";
      POnames[30] = "N563";
      POnames[31] = "N565";
      POnames[32] = "N567";
      POnames[33] = "N569";
      POnames[34] = "N571";
      POnames[35] = "N573";
      POnames[36] = "N582";
      POnames[37] = "N643";
      POnames[38] = "N707";
      POnames[39] = "N813";
      POnames[40] = "N881";
      POnames[41] = "N882";
      POnames[42] = "N883";
      POnames[43] = "N884";
      POnames[44] = "N885";
      POnames[45] = "N889";
      POnames[46] = "N945";
      POnames[47] = "N1110";
      POnames[48] = "N1111";
      POnames[49] = "N1112";
      POnames[50] = "N1113";
      POnames[51] = "N1114";
      POnames[52] = "N1489";
      POnames[53] = "N1490";
      POnames[54] = "N1781";
      POnames[55] = "N10025";
      POnames[56] = "N10101";
      POnames[57] = "N10102";
      POnames[58] = "N10103";
      POnames[59] = "N10104";
      POnames[60] = "N10109";
      POnames[61] = "N10110";
      POnames[62] = "N10111";
      POnames[63] = "N10112";
      POnames[64] = "N10350";
      POnames[65] = "N10351";
      POnames[66] = "N10352";
      POnames[67] = "N10353";
      POnames[68] = "N10574";
      POnames[69] = "N10575";
      POnames[70] = "N10576";
      POnames[71] = "N10628";
      POnames[72] = "N10632";
      POnames[73] = "N10641";
      POnames[74] = "N10704";
      POnames[75] = "N10706";
      POnames[76] = "N10711";
      POnames[77] = "N10712";
      POnames[78] = "N10713";
      POnames[79] = "N10714";
      POnames[80] = "N10715";
      POnames[81] = "N10716";
      POnames[82] = "N10717";
      POnames[83] = "N10718";
      POnames[84] = "N10729";
      POnames[85] = "N10759";
      POnames[86] = "N10760";
      POnames[87] = "N10761";
      POnames[88] = "N10762";
      POnames[89] = "N10763";
      POnames[90] = "N10827";
      POnames[91] = "N10837";
      POnames[92] = "N10838";
      POnames[93] = "N10839";
      POnames[94] = "N10840";
      POnames[95] = "N10868";
      POnames[96] = "N10869";
      POnames[97] = "N10870";
      POnames[98] = "N10871";
      POnames[99] = "N10905";
      POnames[100] = "N10906";
      POnames[101] = "N10907";
      POnames[102] = "N10908";
      POnames[103] = "N11333";
      POnames[104] = "N11334";
      POnames[105] = "N11340";
      POnames[106] = "N11342";
      POnames[107] = "N241_O";
      nofails = 0; pattern = -1; lastpattern = 0;
      prev_pat = -2; error_banner = -2;
      /*** No test setup procedure ***/


      /*** Non-scan test ***/

      if (verbose >= 1) $display("// %t : Begin patterns, first pattern = 0", $time);
pattern = 0; // 0
ALLPIS = 207'b111001010001111110010100101000100111100010000100001101001010001100100101010100111101001110001111100001101001100000101011001010111010101101001010110001111011000000110100001001101101101010001001011101111111111;
XPCT = 108'b110001001110110101000100101101111111100110111111111111101111110000011111100100011010111110011000011101100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 200

pattern = 1; // 200
ALLPIS = 207'b111100101000111111001010010100010011110001000010000110100101000110010010101010011110100111000111110000110100110000010101100101011101010110100101011000111101100000011010000100110110110101000100101110111111111;
XPCT = 108'b111000101011011010100010010110111111101111111101111111000000010110101110110010011111100100111001010010011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 400

pattern = 2; // 400
ALLPIS = 207'b100111000101100001110001100010101110011010100101001110011000101111101100000001110010011101101100011001110011111000100001111000010100000110011000011101100101110000111001001011110110110000101011001010100000000;
XPCT = 108'b110001011011011000010101100110100000011001111100001011111111101000111111111110110000110011111111000000110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 600

pattern = 3; // 600
ALLPIS = 207'b101010110011001110101100011001110000101111010110101010000110011011010011010100000100000000111001101101010000011100111011110110110000101110000110111111001001111000101000101100010110110010011100111000101111111;
XPCT = 108'b110101100011011001001110011100101111001011111100001011001111000001110101011100110110111100011001001111011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 800

pattern = 4; // 800
ALLPIS = 207'b001100001000011001000010100100011111110101101111011000001001000001001100111110111111001110010011010111000001101110110110110001100010111010001001101110011111111100100000011111100110110011000111000001101000000;
XPCT = 108'b000011111011011001100011100001101000100001111001111110000000100011010100010011110011101100111110100111110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1000

pattern = 5; // 1000
ALLPIS = 207'b000110000100001100100001010010001111111010110111101100000100100000100110011111011111100111001001101011100000110111011011011000110001011101000100110111001111111110010000001111110011011001100011100000110100000;
XPCT = 108'b000001111001101100110001110000110100001001011001011010001111111000000101111111000111111000000001101001111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1200

pattern = 6; // 1200
ALLPIS = 207'b111010010011111000000100000001100000011111011111111011001000011100110110011011010010111101101011010100011001111011000110100110100010000011101000101010011100111111111100001110010100000110111000101101100101111;
XPCT = 108'b110001110010000011011100010101100101001110111111011011111111001100000101010101100101110111000001001111100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1400

pattern = 7; // 1400
ALLPIS = 207'b111101001001111100000010000000110000001111101111111101100100001110011011001101101001011110110101101010001100111101100011010011010001000001110100010101001110011111111110000111001010000011011100010110110010111;
XPCT = 108'b111000110101000001101110001010110010100111111111111111100110000100011101011011001101101111111110111110011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1600

pattern = 8; // 1600
ALLPIS = 207'b000111110101000000010101101000111111100101110011110011111000001011101000110010001001100001010101010100101111111110011010100011010010001101110000111011011100001111001011001010001000101011100111010110100110100;
XPCT = 108'b001001010100010101110011101010100110010101101010001010001111011001011011111101111100110011011000101110111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1800

pattern = 9; // 1800
ALLPIS = 207'b100011111010100000001010110100011111110010111001111001111100000101110100011001000100110000101010101010010111111111001101010001101001000110111000011101101110000111100101100101000100010101110011101011010011010;
XPCT = 108'b110100100010001010111001110111010011010011101111010001010110001100011111001000100111101010111110010010100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2000

pattern = 10; // 2000
ALLPIS = 207'b110001111101010000000101011010001111111001011100111100111110000010111010001100100010011000010101010101001011111111100110101000110100100011011100001110110111000011110010110010100010001010111001110101101001101;
XPCT = 108'b111110011001000101011100111001101001100111110101111111101111110011011111001111101000111101111110111011110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2200

pattern = 11; // 2200
ALLPIS = 207'b100001101111010110010110000101100000011110101010010011010101001101111000010010101100000010000101001011001100011111011000011110100000111100100100110110100000100001001101010000111100101111010101100111001011001;
XPCT = 108'b110010001110010111101010110011001011111101111110100101011111011010111111011110001011111101011000010011010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2400

pattern = 12; // 2400
ALLPIS = 207'b001001100110010101011111101010010111101101010001000100100000101010011001011101101011001111001101000100001111101111000111000101101010110011011000101010101011010000010010100001110011111101100011101110011010011;
XPCT = 108'b001100001001111110110001110110011010101111111001111110011001111001011110101111101100110110000000001110111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2600

pattern = 13; // 2600
ALLPIS = 207'b100100110011001010101111110101001011110110101000100010010000010101001100101110110101100111100110100010000111110111100011100010110101011001101100010101010101101000001001010000111001111110110001110111001101001;
XPCT = 108'b110010001100111111011000111011001101111111001100101111011111101001111111101100111011110000111110100111000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2800

pattern = 14; // 2800
ALLPIS = 207'b101011001000011011000011010010000010011001010000011100000010000110000011000011100111111101111100110000101010011011011010111011100000000001111100111011010001110100110000100001110001010101010001100110011001011;
XPCT = 108'b110100001000101010101000110010011001001101111101011011111001000100011110001111100110110011000000010101001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3000

pattern = 15; // 3000
ALLPIS = 207'b110101100100001101100001101001000001001100101000001110000001000011000001100001110011111110111110011000010101001101101101011101110000000000111110011101101000111010011000010000111000101010101000110011001100101;
XPCT = 108'b110010001100010101010100011011001100101011111101111111100110010101111111101000011111100010011111010011001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3200

pattern = 16; // 3200
ALLPIS = 207'b000011100011111000100100011100000111000100010000001010001010101101000101100100000100110001010000101101100011000110011101100100000010101101010101111111001111011101111000000001110001111111011101000100011001101;
XPCT = 108'b000000001000111111101110100000011001001101111000001010001111111110101111001110110101110000111110110111001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3400

pattern = 17; // 3400
ALLPIS = 207'b011000100000000010000110100110100100000000001100001000001111011010000111100110111111010110100111110111011000000011100101111000111011111011100000001110011100101110001000001001010101010101100111111111110011001;
XPCT = 108'b000001000010101010110011111111110011101111111001111110001111101000101111110100000111110101100000101001101001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3600

pattern = 18; // 3600
ALLPIS = 207'b001100010000000001000011010011010010000000000110000100000111101101000011110011011111101011010011111011101100000001110010111100011101111101110000000111001110010111000100000100101010101010110011111111111001100;
XPCT = 108'b000000101101010101011001111111111001100101111001111110000000111111011110011011011111101010011110100111000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3800

pattern = 19; // 3800
ALLPIS = 207'b100110001000000000100001101001101001000000000011000010000011110110100001111001101111110101101001111101110110000000111001011110001110111110111000000011100111001011100010000010010101010101011001111111111100110;
XPCT = 108'b111000010010101010101100111111111100001101111101011011010000001010001110010000001111100101111000000010011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4000

pattern = 20; // 4000
ALLPIS = 207'b010011000100000000010000110100110100100000000001100001000001111011010000111100110111111010110100111110111011000000011100101111000111011111011100000001110011100101110001000001001010101010101100111111111110011;
XPCT = 108'b000000000101010101010110011111111110010110111011011010011001011100011110000100101010111110000000010100011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4200

pattern = 21; // 4200
ALLPIS = 207'b101001100010000000001000011010011010010000000000110000100000111101101000011110011011111101011010011111011101100000001110010111100011101111101110000000111001110010111000100000100101010101010110011111111111001;
XPCT = 108'b110100001010101010101011001111111111100110111100101111111111011111011111000100011101111111100000000100000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4400

pattern = 22; // 4400
ALLPIS = 207'b001101100000111110010000100101101010101010000100010101011010010010010001011011110000110000100010101110000111010000101100000001001011011010111101110001100111111001101000011001111111000000100010010010000000011;
XPCT = 108'b000011001111100000010001001010000000101001111010101110010000011101101110011000010001101111111110000011101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4600

pattern = 23; // 4600
ALLPIS = 207'b011111100001100001011100111010010010110111000110000111100111000101101101111001000101010110011110110110101010001000111101001010011111000000010100001001001000111100000000000101010010001010011000010100111111110;
XPCT = 108'b000000100001000101001100001000111111001111111011011010001111011010111111110100001101111100000111100000000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4800

pattern = 24; // 4800
ALLPIS = 207'b110110100001001110111010110101101110111001100111001110111001101110010011101000011111100101000000111010111100100100110101101111110101001101000000110101011111011110110100001011000100101111000101010111100000000;
XPCT = 108'b110001010010010111100010101011100000000111111101011011001111001101001111111110000111110010111110101110001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5000

pattern = 25; // 5000
ALLPIS = 207'b011011010000100111011101011010110111011100110011100111011100110111001001110100001111110010100000011101011110010010011010110111111010100110100000011010101111101111011010000101100010010111100010101011110000000;
XPCT = 108'b001000101001001011110001010111110000000011111011011010011111110110011111001110111000110110000001011000000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5200

pattern = 26; // 5200
ALLPIS = 207'b110100111001101101111010000101111100001100011101111110100100010111000001101110111010110111011111101111000110101001100110010001000111111110011010111100101100110111011001001011011100100001111000001000000111111;
XPCT = 108'b110001010110010000111100000100000111111011111101111111001111100011111011100101100111111110100111011111011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5400

pattern = 27; // 5400
ALLPIS = 207'b011010011100110110111101000010111110000110001110111111010010001011100000110111011101011011101111110111100011010100110011001000100011111111001101011110010110011011101100100101101110010000111100000100000011111;
XPCT = 108'b000100101111001000011110000000000011000111010011011010010110110010101111010000011100101101111110110101010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5600

pattern = 28; // 5600
ALLPIS = 207'b010100011111100101001010001001111000100001000011010010100011001001010101001111010011100011111000011010011000001010110010101110101011010010101100011110110000001101000010011011011010100010010111011111111110000;
XPCT = 108'b001011010101010001001011101111111110101111111001111110001111000101101111110101010011111110011110110011110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5800

pattern = 29; // 5800
ALLPIS = 207'b001010001111110010100101000100111100010000100001101001010001100100101010100111101001110001111100001101001100000101011001010111010101101001010110001111011000000110100001001101101101010001001011101111111111000;
XPCT = 108'b000001101110101000100101110111111111010101111011011010011111110011001111000100010101111101011110001001111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6000

pattern = 30; // 6000
ALLPIS = 207'b100101000111111001010010100010011110001000010000110100101000110010010101010011110100111000111110000110100110000010101100101011101010110100101011000111101100000011010000100110110110101000100101110111111111100;
XPCT = 108'b110100111011010100010010111011111111101101111101111111101111101000011111010111010001111001111110111110001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6200

pattern = 31; // 6200
ALLPIS = 207'b110010100011111100101001010001001111000100001000011010010100011001001010101001111010011100011111000011010011000001010110010101110101011010010101100011110110000001101000010011011011010100010010111011111111110;
XPCT = 108'b110010010101101010001001011111111111001011111101011011111111101001001111111111101011110100000110000111000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6400

pattern = 32; // 6400
ALLPIS = 207'b000011001000000000001010010010000111011011010010001010000100110011010110001110000011110100101001001000011100000000110011110010000010001001100001100111111011110000001000100000110101010100100011000001101100010;
XPCT = 108'b000100001010101010010001100001101100001011111000001010011001111010111100010110010100111101000000001001101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6600

pattern = 33; // 6600
ALLPIS = 207'b100001100100000000000101001001000011101101101001000101000010011001101011000111000001111010010100100100001110000000011001111001000001000100110000110011111101111000000100010000011010101010010001100000110110001;
XPCT = 108'b110010000101010101001000110000110110101001111111111111110000010100011110000010111101100110011110111110000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6800

pattern = 34; // 6800
ALLPIS = 207'b110011111010000000001000110110100110101101100110101000100101111111100011101101100011001001100011011010011011000000111111001110100010101011111001111110000101001100001010101000111000000001101011110001110111010;
XPCT = 108'b111101001100000000110101111001110111001011111101011011111001011001011110110100010110110110000000000100110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7000

pattern = 35; // 7000
ALLPIS = 207'b011010110101000000001110001001010100001101100001011110010110001100100111111000110010010000011000100101010001100000101100010101010011011100011101011000111001010110001101110100101001010100010110111001010111111;
XPCT = 108'b000110101100101010001011011101010111010011111001011010001111010011110101000100101010110101111001100101100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7200

pattern = 36; // 7200
ALLPIS = 207'b101110010010100000001101010110101101011101100010100101001111110101000101110010011010111100100101011010110100110000100101111000101011100111101111001011100111011011001110011010100001111110101000011101000111101;
XPCT = 108'b111011011000111111010100001101000111000111111110001011110000110101000100010010110001100000011111110001001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7400

pattern = 37; // 7400
ALLPIS = 207'b010111001001010000000110101011010110101110110001010010100111111010100010111001001101011110010010101101011010011000010010111100010101110011110111100101110011101101100111001101010000111111010100001110100011110;
XPCT = 108'b001001100000011111101010000110100011011111111001011010001111001111101111010111010110110101111001111000101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7600

pattern = 38; // 7600
ALLPIS = 207'b100100010110010100000100100011110110000110000101010001101011100111000011101001010010101101110000001111011000100110011101010110000100011000001101001010100001000011011101100011001110100101100100100011011110110;
XPCT = 108'b110100010111010010110010010011011110110001111110101111110110100000101111101000111100100110011000111011100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7800

pattern = 39; // 7800
ALLPIS = 207'b011000100001100101000100000001111110001100001000010001011000100000011011111101010101010001001000100111111000001001111110101100100000000010110011100001010101101000110011001000101001000011001000101000000001100;
XPCT = 108'b001001001100100001100100010100000001110011111011111110001111000011001111100101010101111111111110001010001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8000

pattern = 40; // 8000
ALLPIS = 207'b001100010000110010100010000000111111000110000100001000101100010000001101111110101010101000100100010011111100000100111111010110010000000001011001110000101010110100011001100100010100100001100100010100000000110;
XPCT = 108'b000100100010010000110010001000000000111101111000101110000000100101111110000001011110101111111000000000011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8200

pattern = 41; // 8200
ALLPIS = 207'b100101000000011001011011010010011000111000010000001110010010111011010000110001010110100000111011000001100010000010101100011001001010001001001101011111101110101010000100010010111111000100010001001011101100001;
XPCT = 108'b110010011111100010001000100111101100101011111101111111010110011110001111111001101111101100111111000001000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8400

pattern = 42; // 8400
ALLPIS = 207'b110001101000001100100111111011001011000111011010001101001101101110111110010110101000100100110100101000101101000001100101111110100111001101000111001000001100100101001010101001101010110110101011100100011010010;
XPCT = 108'b111101001101011011010101110000011010100111111111111111010000111110101110011000111000101111011111111011011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8600

pattern = 43; // 8600
ALLPIS = 207'b111000110100000110010011111101100101100011101101000110100110110111011111001011010100010010011010010100010110100000110010111111010011100110100011100100000110010010100101010100110101011011010101110010001101001;
XPCT = 108'b110010101010101101101010111010001101111011111101111111001111001100010101101101001011111001100001111001010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8800

pattern = 44; // 8800
ALLPIS = 207'b111111010010000011000011101100110101101010100100101001010111101000111001101011101001111101100100000010010111010000101010101101101011111010110000010101111000111001011010001010101111111001001001111000101010110;
XPCT = 108'b111001011111111100100100111100101010000011111111011011100000010101011110010000100101101000100110000110011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9000

pattern = 45; // 9000
ALLPIS = 207'b111100111100100000111010101001001010000001111011000000010001001001011000010100111001101011110000001000111001110100111001011001011000110111001101100010100101111110011110000010011110101010110001011111100110111;
XPCT = 108'b111000010111010101011000101111100110101111011101111111110000010001110100110011001111101010000111100001101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9200

pattern = 46; // 9200
ALLPIS = 207'b111101010110010000010111000110100010011011101111101010001100010111111010000100011111000001010001001100000000111010101111011110101110010010000111010110101001001111000111100001111010000001111011101110011111001;
XPCT = 108'b111100001101000000111101110110011111111111111101111111010000011111011110010000011110100000011111100110101001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9400

pattern = 47; // 9400
ALLPIS = 207'b111110101011001000001011100011010001001101110111110101000110001011111101000010001111100000101000100110000000011101010111101111010111001001000011101011010100100111100011110000111101000000111101110111001111100;
XPCT = 108'b111110001110100000011110111011001111011111111111011011001111011011000101001110111000111111011001010101001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9600

pattern = 48; // 9600
ALLPIS = 207'b011111010101100100000101110001101000100110111011111010100011000101111110100001000111110000010100010011000000001110101011110111101011100100100001110101101010010011110001111000011110100000011110111011100111110;
XPCT = 108'b000111000111010000001111011111100111011011111001011010001001010110111110000111110010111110111001101100001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9800

pattern = 49; // 9800
ALLPIS = 207'b001111101010110010000010111000110100010011011101111101010001100010111111010000100011111000001010001001100000000111010101111011110101110010010000111010110101001001111000111100001111010000001111011101110011111;
XPCT = 108'b000111100111101000000111101101110011000101111010000000000000110110001010111000110000101101011001011011011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10000

pattern = 50; // 10000
ALLPIS = 207'b100111110101011001000001011100011010001001101110111110101000110001011111101000010001111100000101000100110000000011101010111101111010111001001000011101011010100100111100011110000111101000000111101110111001111;
XPCT = 108'b110011110011110100000011110110111001000101111100001011100110110000101111001000111000101011011110000100000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10200

pattern = 51; // 10200
ALLPIS = 207'b110000110010101100101010111100001010011111100101010101010000101011111001111010001011001010101011101010000100000001000110101100111111010101000101101001010110100010010110101111110110100000100000110110110000101;
XPCT = 108'b111101111011010000010000011010110000101111111111111111111111010111111111011110000100111110000000000010111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10400

pattern = 52; // 10400
ALLPIS = 207'b111011010001010110011111001100000010010100100000100000101100100110101010110011000110010001111100111101011110000000010000100100011101100011000011010011010000100001000011110111001110000100110011011010110100000;
XPCT = 108'b111110110111000010011001101110110100010011111101011011011111110101101111000111110111110011111110101101010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10600

pattern = 53; // 10600
ALLPIS = 207'b011110100000101011000101110100000110010001000010011010010010100000000011010111100000111100010111010110110011000000111011100000001100111000000000001110010011100000101001011011010010010110111010101100110110010;
XPCT = 108'b000011010001001011011101010100110110011111111001011010000000010110111110000011010011100101000111110100100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10800

pattern = 54; // 10800
ALLPIS = 207'b001111010000010101100010111010000011001000100001001101001001010000000001101011110000011110001011101011011001100000011101110000000110011100000000000111001001110000010100101101101001001011011101010110011011001;
XPCT = 108'b000101101100100101101110101010011011000101111011011010010000000111001110010001110100101011011111101001011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11000

pattern = 55; // 11000
ALLPIS = 207'b000100100000001010111011001111000110111111000010101100100000011011010110111011111011111011101100111101110000110000111101001010000001000111100001100100011111001000000010110110000001110001001101101010100001110;
XPCT = 108'b001110110000111000100110110110100001100011111001111110010000011101001010110000011010101100100111000000011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11200

pattern = 56; // 11200
ALLPIS = 207'b100010010000000101011101100111100011011111100001010110010000001101101011011101111101111101110110011110111000011000011110100101000000100011110000110010001111100100000001011011000000111000100110110101010000111;
XPCT = 108'b110011010000011100010011011001010000010111111101011011100000000100001110001011100011101000111001011101110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11400

pattern = 57; // 11400
ALLPIS = 207'b011001000000000001010010010000111011011010010001010000100110011010110001110000011110100101001001000011100000000110011110010000010001001100001100111111011110000001000100000110101010100100011000001101100010000;
XPCT = 108'b000000111101010010001100000101100010100111111001111110010110101001111101111010001111101000011111001111100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11600

pattern = 58; // 11600
ALLPIS = 207'b000110010000000000010100100100001110110110100100010100001001100110101100011100000111101001010010010000111000000001100111100100000100010011000011001111110111100000010001000001101010101001000110000011011000100;
XPCT = 108'b000000001101010100100011000011011000010001111001011010011111100111001111100101111111111010000000111111011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11800

pattern = 59; // 11800
ALLPIS = 207'b000110111011011010110011101001001010100111100000110011110000010100101111011010111110101100011100011010100111010110101010110111000000100000010011110001101101010111100101111111110011000001000000011000110101000;
XPCT = 108'b000111111001100000100000001100110101011001111011011010001111111011001111001100100000111111011111110111001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12000

pattern = 60; // 12000
ALLPIS = 207'b000011011101101101011001110100100101010011110000011001111000001010010111101101011111010110001110001101010011101011010101011011100000010000001001111000110110101011110010111111111001100000100000001100011010100;
XPCT = 108'b001111111100110000010000000100011010001111111011011010001111101010101011001101100001110100011000000001001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12200

pattern = 61; // 12200
ALLPIS = 207'b100111010101101100011111010011011000001110011000111111001100010001100100101100010001000111011011011100001110100011000000011010110000101000010111001101110110000010011100100000001111110001010000011110111000010;
XPCT = 108'b110100000111111000101000001110111000000111111110001011011111111111111111101100101110111101011001111101001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12400

pattern = 62; // 12400
ALLPIS = 207'b010101010001101100111100000000100110100000101100101100010110011100011101001100110110001111110001110100100000000111001010111010011000110100011000010111010110010110101011101111110100111001101000010111101001001;
XPCT = 108'b001101111010011100110100001011101001111111111001111110011111000000010111111100110111111100011000000100000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12600

pattern = 63; // 12600
ALLPIS = 207'b110110001001110110010110110100101100111011111011010010111101101101010000111110010010110101110010010000011011101010100111110101000110011101001111111101000011001110011000000100000100101110111010001001100000110;
XPCT = 108'b110000100010010111011101000101100000000011111101011011011111001001001111111101101111110010011000000010011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12800

pattern = 64; // 12800
ALLPIS = 207'b101110111111110000111100011001101110011101001110101101010111010001000011100010111011111011010010101001010101010001111100100110110001110111011010000111100110011000010100111110111000101011001110101110000010101;
XPCT = 108'b110111111100010101100111010110000010001111111111011011101111101100110101011100010000111011011000000011111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13000

pattern = 65; // 13000
ALLPIS = 207'b010001100100100010101101100101111101101001000111100101011011111100001110101011100011010001110101001110001101111110010100100100011000011011111110110010011110011011101111100000101111010100100111001111110100010;
XPCT = 108'b001100001111101010010011100111110100110111111011111110011001000101101110111101001011110011000000011100011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13200

pattern = 66; // 13200
ALLPIS = 207'b101000110010010001010110110010111110110100100011110010101101111110000111010101110001101000111010100111000110111111001010010010001100001101111111011001001111001101110111110000010111101010010011100111111010001;
XPCT = 108'b111110000011110101001001110011111010111101101101111111111111101111111111000111001010111001100000110101111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13400

pattern = 67; // 13400
ALLPIS = 207'b010000010000010010110000010101111100000001011010011010001110111000100100000110100111111011101010100001100110000101000011011111011000101000111010111001001001000010111100111111000100001110011001000100001000011;
XPCT = 108'b000111110010000111001100100000001000100111111001111110010110001111101111011001110010100011100110110011100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13600

pattern = 68; // 13600
ALLPIS = 207'b101110110011010011101011100011110100100111001101111110110111001000111101011001101101010001101001001010010100010100001011011000101100110100001110101101001001110110111011100000010001000110001100111010110001001;
XPCT = 108'b111100000000100011000110011110110001011011110100000001011111000111000101101111101110110111111001001000001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13800

pattern = 69; // 13800
ALLPIS = 207'b011100000100001011011101110000011100010100001010010001011111101001111111110111001011000100000111110111101001100111110111101101111001010101101110111111001100101100101000000111000010001010010100011100111110011;
XPCT = 108'b000000110001000101001010001100111110100111011011111110010000010110000100011000111101101100000000001101111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14000

pattern = 70; // 14000
ALLPIS = 207'b001110000010000101101110111000001110001010000101001000101111110100111111111011100101100010000011111011110100110011111011110110111100101010110111011111100110010110010100000011100001000101001010001110011111001;
XPCT = 108'b000000011000100010100101000110011111000111111001010000000000101100100100011011111111100111011111000010100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14200

pattern = 71; // 14200
ALLPIS = 207'b110101011011111011101000000111001001000101000001100001111011101001100000100100000111110100111100100100011010011010010100001010101111101010111110000110010100110010000000111111001011010000010010111011010010110;
XPCT = 108'b110111110101101000001001011111010010100011111111111111000110000001101111001010101100101101011111011001101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14400

pattern = 72; // 14400
ALLPIS = 207'b100000110111011000100111101110001101111110110000111111010101111101100111010101010110101101101011001101001011110000011100011100100010010010111110101011100010111011101000001100001101000100011001010110010011110;
XPCT = 108'b110001100110100010001100101010010011100101111110101111101111100000111111110111110101110110011000110011101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14600

pattern = 73; // 14600
ALLPIS = 207'b010000011011101100010011110111000110111111011000011111101010111110110011101010101011010110110101100110100101111000001110001110010001001001011111010101110001011101110100000110000110100010001100101011001001111;
XPCT = 108'b000000110011010001000110010111001001100011111011111110011111111110011111111101001101111110100001100010001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14800

pattern = 74; // 14800
ALLPIS = 207'b101110110110101100111010010010101001111000001100111100000101001011110110101111101011000111000110101001110101101010101101110000001000000100111100011011010101111001011111111100110000010000000110001101010001111;
XPCT = 108'b111111101000001000000011000101010001011111111100000001010000111010011010101000000010101110111000100111111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15000

pattern = 75; // 15000
ALLPIS = 207'b011011101101101011001110100100101010011110000011001111000001010010111101101011111010110001110001101010011101011010101011011100000010000001001111000110110101011110010111111111001100000100000001100011010100011;
XPCT = 108'b001111110110000010000000110011010100010011111011011010010110110111111111111001110100100111011111011100101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15200

pattern = 76; // 15200
ALLPIS = 207'b001101110110110101100111010010010101001111000001100111100000101001011110110101111101011000111000110101001110101101010101101110000001000000100111100011011010101111001011111111100110000010000000110001101010001;
XPCT = 108'b001111111011000001000000011001101010110001111010101110010000111011101110000011110000101111111111100100011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15400

      $display("// %t : Simulation of %0d patterns completed with %0d errors\n", $time, pattern+1, nofails);
      if (verbose >=2) $finish(2);
      /* else */ $finish(0);
   end
endmodule
