// Verilog pattern output written by  TetraMAX (TM)  B-2008.09-SP2-i081128_181834 
// Date: Wed Jul  6 12:11:51 2011
// Module tested: c7552

//     Uncollapsed Stuck Fault Summary Report
// -----------------------------------------------
// fault class                     code   #faults
// ------------------------------  ----  ---------
// Detected                         DT       6858
// Possibly detected                PT          0
// Undetectable                     UD          0
// ATPG untestable                  AU          0
// Not detected                     ND         30
// -----------------------------------------------
// total faults                              6888
// test coverage                            99.56%
// -----------------------------------------------
// 
//            Pattern Summary Report
// -----------------------------------------------
// #internal patterns                         259
//     #basic_scan patterns                   259
// -----------------------------------------------
// 
// There are no rule fails
// There are no clocks
// There are no constraint ports
// There are no equivalent pins
// There are no net connections

`timescale 1 ns / 1 ns

//
// --- NOTE: Remove the comment to define 'tmax_iddq' to activate processing of IDDQ events
//     Or use '+define+tmax_iddq' on the verilog compile line
//
//`define tmax_iddq

module AAA_tmax_testbench_1_16 ;
   parameter NAMELENGTH = 200; // max length of names reported in fails
   integer nofails, bit, pattern, lastpattern;
   integer error_banner; // flag for tracking displayed error banner
   integer loads;        // number of load_unloads for current pattern
   integer patm1;        // pattern - 1
   integer patp1;        // pattern + lastpattern
   integer prev_pat;     // previous pattern number
   integer report_interval; // report pattern progress every Nth pattern
   integer verbose;      // message verbosity level
   parameter NINPUTS = 207, NOUTPUTS = 108;
   wire [0:NOUTPUTS-1] PO; reg [0:NOUTPUTS-1] ALLPOS, XPCT, MASK;
   reg [0:NINPUTS-1] PI, ALLPIS;
   reg [0:8*(NAMELENGTH-1)] POnames [0:NOUTPUTS-1];
   event IDDQ;

   wire N1;
   wire N5;
   wire N9;
   wire N12;
   wire N15;
   wire N18;
   wire N23;
   wire N26;
   wire N29;
   wire N32;
   wire N35;
   wire N38;
   wire N41;
   wire N44;
   wire N47;
   wire N50;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N69;
   wire N70;
   wire N73;
   wire N74;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N82;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N94;
   wire N97;
   wire N100;
   wire N103;
   wire N106;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N118;
   wire N121;
   wire N124;
   wire N127;
   wire N130;
   wire N133;
   wire N134;
   wire N135;
   wire N138;
   wire N141;
   wire N144;
   wire N147;
   wire N150;
   wire N151;
   wire N152;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N178;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire N185;
   wire N186;
   wire N187;
   wire N188;
   wire N189;
   wire N190;
   wire N191;
   wire N192;
   wire N193;
   wire N194;
   wire N195;
   wire N196;
   wire N197;
   wire N198;
   wire N199;
   wire N200;
   wire N201;
   wire N202;
   wire N203;
   wire N204;
   wire N205;
   wire N206;
   wire N207;
   wire N208;
   wire N209;
   wire N210;
   wire N211;
   wire N212;
   wire N213;
   wire N214;
   wire N215;
   wire N216;
   wire N217;
   wire N218;
   wire N219;
   wire N220;
   wire N221;
   wire N222;
   wire N223;
   wire N224;
   wire N225;
   wire N226;
   wire N227;
   wire N228;
   wire N229;
   wire N230;
   wire N231;
   wire N232;
   wire N233;
   wire N234;
   wire N235;
   wire N236;
   wire N237;
   wire N238;
   wire N239;
   wire N240;
   wire N242;
   wire N245;
   wire N248;
   wire N251;
   wire N254;
   wire N257;
   wire N260;
   wire N263;
   wire N267;
   wire N271;
   wire N274;
   wire N277;
   wire N280;
   wire N283;
   wire N286;
   wire N289;
   wire N293;
   wire N296;
   wire N299;
   wire N303;
   wire N307;
   wire N310;
   wire N313;
   wire N316;
   wire N319;
   wire N322;
   wire N325;
   wire N328;
   wire N331;
   wire N334;
   wire N337;
   wire N340;
   wire N343;
   wire N346;
   wire N349;
   wire N352;
   wire N355;
   wire N358;
   wire N361;
   wire N364;
   wire N367;
   wire N382;
   wire N241_I;
   wire N387;
   wire N388;
   wire N478;
   wire N482;
   wire N484;
   wire N486;
   wire N489;
   wire N492;
   wire N501;
   wire N505;
   wire N507;
   wire N509;
   wire N511;
   wire N513;
   wire N515;
   wire N517;
   wire N519;
   wire N535;
   wire N537;
   wire N539;
   wire N541;
   wire N543;
   wire N545;
   wire N547;
   wire N549;
   wire N551;
   wire N553;
   wire N556;
   wire N559;
   wire N561;
   wire N563;
   wire N565;
   wire N567;
   wire N569;
   wire N571;
   wire N573;
   wire N582;
   wire N643;
   wire N707;
   wire N813;
   wire N881;
   wire N882;
   wire N883;
   wire N884;
   wire N885;
   wire N889;
   wire N945;
   wire N1110;
   wire N1111;
   wire N1112;
   wire N1113;
   wire N1114;
   wire N1489;
   wire N1490;
   wire N1781;
   wire N10025;
   wire N10101;
   wire N10102;
   wire N10103;
   wire N10104;
   wire N10109;
   wire N10110;
   wire N10111;
   wire N10112;
   wire N10350;
   wire N10351;
   wire N10352;
   wire N10353;
   wire N10574;
   wire N10575;
   wire N10576;
   wire N10628;
   wire N10632;
   wire N10641;
   wire N10704;
   wire N10706;
   wire N10711;
   wire N10712;
   wire N10713;
   wire N10714;
   wire N10715;
   wire N10716;
   wire N10717;
   wire N10718;
   wire N10729;
   wire N10759;
   wire N10760;
   wire N10761;
   wire N10762;
   wire N10763;
   wire N10827;
   wire N10837;
   wire N10838;
   wire N10839;
   wire N10840;
   wire N10868;
   wire N10869;
   wire N10870;
   wire N10871;
   wire N10905;
   wire N10906;
   wire N10907;
   wire N10908;
   wire N11333;
   wire N11334;
   wire N11340;
   wire N11342;
   wire N241_O;

   // map PI[] vector to DUT inputs and bidis
   assign N1 = PI[0];
   assign N5 = PI[1];
   assign N9 = PI[2];
   assign N12 = PI[3];
   assign N15 = PI[4];
   assign N18 = PI[5];
   assign N23 = PI[6];
   assign N26 = PI[7];
   assign N29 = PI[8];
   assign N32 = PI[9];
   assign N35 = PI[10];
   assign N38 = PI[11];
   assign N41 = PI[12];
   assign N44 = PI[13];
   assign N47 = PI[14];
   assign N50 = PI[15];
   assign N53 = PI[16];
   assign N54 = PI[17];
   assign N55 = PI[18];
   assign N56 = PI[19];
   assign N57 = PI[20];
   assign N58 = PI[21];
   assign N59 = PI[22];
   assign N60 = PI[23];
   assign N61 = PI[24];
   assign N62 = PI[25];
   assign N63 = PI[26];
   assign N64 = PI[27];
   assign N65 = PI[28];
   assign N66 = PI[29];
   assign N69 = PI[30];
   assign N70 = PI[31];
   assign N73 = PI[32];
   assign N74 = PI[33];
   assign N75 = PI[34];
   assign N76 = PI[35];
   assign N77 = PI[36];
   assign N78 = PI[37];
   assign N79 = PI[38];
   assign N80 = PI[39];
   assign N81 = PI[40];
   assign N82 = PI[41];
   assign N83 = PI[42];
   assign N84 = PI[43];
   assign N85 = PI[44];
   assign N86 = PI[45];
   assign N87 = PI[46];
   assign N88 = PI[47];
   assign N89 = PI[48];
   assign N94 = PI[49];
   assign N97 = PI[50];
   assign N100 = PI[51];
   assign N103 = PI[52];
   assign N106 = PI[53];
   assign N109 = PI[54];
   assign N110 = PI[55];
   assign N111 = PI[56];
   assign N112 = PI[57];
   assign N113 = PI[58];
   assign N114 = PI[59];
   assign N115 = PI[60];
   assign N118 = PI[61];
   assign N121 = PI[62];
   assign N124 = PI[63];
   assign N127 = PI[64];
   assign N130 = PI[65];
   assign N133 = PI[66];
   assign N134 = PI[67];
   assign N135 = PI[68];
   assign N138 = PI[69];
   assign N141 = PI[70];
   assign N144 = PI[71];
   assign N147 = PI[72];
   assign N150 = PI[73];
   assign N151 = PI[74];
   assign N152 = PI[75];
   assign N153 = PI[76];
   assign N154 = PI[77];
   assign N155 = PI[78];
   assign N156 = PI[79];
   assign N157 = PI[80];
   assign N158 = PI[81];
   assign N159 = PI[82];
   assign N160 = PI[83];
   assign N161 = PI[84];
   assign N162 = PI[85];
   assign N163 = PI[86];
   assign N164 = PI[87];
   assign N165 = PI[88];
   assign N166 = PI[89];
   assign N167 = PI[90];
   assign N168 = PI[91];
   assign N169 = PI[92];
   assign N170 = PI[93];
   assign N171 = PI[94];
   assign N172 = PI[95];
   assign N173 = PI[96];
   assign N174 = PI[97];
   assign N175 = PI[98];
   assign N176 = PI[99];
   assign N177 = PI[100];
   assign N178 = PI[101];
   assign N179 = PI[102];
   assign N180 = PI[103];
   assign N181 = PI[104];
   assign N182 = PI[105];
   assign N183 = PI[106];
   assign N184 = PI[107];
   assign N185 = PI[108];
   assign N186 = PI[109];
   assign N187 = PI[110];
   assign N188 = PI[111];
   assign N189 = PI[112];
   assign N190 = PI[113];
   assign N191 = PI[114];
   assign N192 = PI[115];
   assign N193 = PI[116];
   assign N194 = PI[117];
   assign N195 = PI[118];
   assign N196 = PI[119];
   assign N197 = PI[120];
   assign N198 = PI[121];
   assign N199 = PI[122];
   assign N200 = PI[123];
   assign N201 = PI[124];
   assign N202 = PI[125];
   assign N203 = PI[126];
   assign N204 = PI[127];
   assign N205 = PI[128];
   assign N206 = PI[129];
   assign N207 = PI[130];
   assign N208 = PI[131];
   assign N209 = PI[132];
   assign N210 = PI[133];
   assign N211 = PI[134];
   assign N212 = PI[135];
   assign N213 = PI[136];
   assign N214 = PI[137];
   assign N215 = PI[138];
   assign N216 = PI[139];
   assign N217 = PI[140];
   assign N218 = PI[141];
   assign N219 = PI[142];
   assign N220 = PI[143];
   assign N221 = PI[144];
   assign N222 = PI[145];
   assign N223 = PI[146];
   assign N224 = PI[147];
   assign N225 = PI[148];
   assign N226 = PI[149];
   assign N227 = PI[150];
   assign N228 = PI[151];
   assign N229 = PI[152];
   assign N230 = PI[153];
   assign N231 = PI[154];
   assign N232 = PI[155];
   assign N233 = PI[156];
   assign N234 = PI[157];
   assign N235 = PI[158];
   assign N236 = PI[159];
   assign N237 = PI[160];
   assign N238 = PI[161];
   assign N239 = PI[162];
   assign N240 = PI[163];
   assign N242 = PI[164];
   assign N245 = PI[165];
   assign N248 = PI[166];
   assign N251 = PI[167];
   assign N254 = PI[168];
   assign N257 = PI[169];
   assign N260 = PI[170];
   assign N263 = PI[171];
   assign N267 = PI[172];
   assign N271 = PI[173];
   assign N274 = PI[174];
   assign N277 = PI[175];
   assign N280 = PI[176];
   assign N283 = PI[177];
   assign N286 = PI[178];
   assign N289 = PI[179];
   assign N293 = PI[180];
   assign N296 = PI[181];
   assign N299 = PI[182];
   assign N303 = PI[183];
   assign N307 = PI[184];
   assign N310 = PI[185];
   assign N313 = PI[186];
   assign N316 = PI[187];
   assign N319 = PI[188];
   assign N322 = PI[189];
   assign N325 = PI[190];
   assign N328 = PI[191];
   assign N331 = PI[192];
   assign N334 = PI[193];
   assign N337 = PI[194];
   assign N340 = PI[195];
   assign N343 = PI[196];
   assign N346 = PI[197];
   assign N349 = PI[198];
   assign N352 = PI[199];
   assign N355 = PI[200];
   assign N358 = PI[201];
   assign N361 = PI[202];
   assign N364 = PI[203];
   assign N367 = PI[204];
   assign N382 = PI[205];
   assign N241_I = PI[206];

   // map DUT outputs and bidis to PO[] vector
   assign
      PO[0] = N387 ,
      PO[1] = N388 ,
      PO[2] = N478 ,
      PO[3] = N482 ,
      PO[4] = N484 ,
      PO[5] = N486 ,
      PO[6] = N489 ,
      PO[7] = N492 ,
      PO[8] = N501 ,
      PO[9] = N505 ,
      PO[10] = N507 ,
      PO[11] = N509 ,
      PO[12] = N511 ,
      PO[13] = N513 ,
      PO[14] = N515 ,
      PO[15] = N517 ,
      PO[16] = N519 ,
      PO[17] = N535 ,
      PO[18] = N537 ,
      PO[19] = N539 ,
      PO[20] = N541 ,
      PO[21] = N543 ,
      PO[22] = N545 ,
      PO[23] = N547 ,
      PO[24] = N549 ,
      PO[25] = N551 ,
      PO[26] = N553 ,
      PO[27] = N556 ,
      PO[28] = N559 ,
      PO[29] = N561 ,
      PO[30] = N563 ,
      PO[31] = N565 ;
   assign
      PO[32] = N567 ,
      PO[33] = N569 ,
      PO[34] = N571 ,
      PO[35] = N573 ,
      PO[36] = N582 ,
      PO[37] = N643 ,
      PO[38] = N707 ,
      PO[39] = N813 ,
      PO[40] = N881 ,
      PO[41] = N882 ,
      PO[42] = N883 ,
      PO[43] = N884 ,
      PO[44] = N885 ,
      PO[45] = N889 ,
      PO[46] = N945 ,
      PO[47] = N1110 ,
      PO[48] = N1111 ,
      PO[49] = N1112 ,
      PO[50] = N1113 ,
      PO[51] = N1114 ,
      PO[52] = N1489 ,
      PO[53] = N1490 ,
      PO[54] = N1781 ,
      PO[55] = N10025 ,
      PO[56] = N10101 ,
      PO[57] = N10102 ,
      PO[58] = N10103 ,
      PO[59] = N10104 ,
      PO[60] = N10109 ,
      PO[61] = N10110 ,
      PO[62] = N10111 ,
      PO[63] = N10112 ;
   assign
      PO[64] = N10350 ,
      PO[65] = N10351 ,
      PO[66] = N10352 ,
      PO[67] = N10353 ,
      PO[68] = N10574 ,
      PO[69] = N10575 ,
      PO[70] = N10576 ,
      PO[71] = N10628 ,
      PO[72] = N10632 ,
      PO[73] = N10641 ,
      PO[74] = N10704 ,
      PO[75] = N10706 ,
      PO[76] = N10711 ,
      PO[77] = N10712 ,
      PO[78] = N10713 ,
      PO[79] = N10714 ,
      PO[80] = N10715 ,
      PO[81] = N10716 ,
      PO[82] = N10717 ,
      PO[83] = N10718 ,
      PO[84] = N10729 ,
      PO[85] = N10759 ,
      PO[86] = N10760 ,
      PO[87] = N10761 ,
      PO[88] = N10762 ,
      PO[89] = N10763 ,
      PO[90] = N10827 ,
      PO[91] = N10837 ,
      PO[92] = N10838 ,
      PO[93] = N10839 ,
      PO[94] = N10840 ,
      PO[95] = N10868 ;
   assign
      PO[96] = N10869 ,
      PO[97] = N10870 ,
      PO[98] = N10871 ,
      PO[99] = N10905 ,
      PO[100] = N10906 ,
      PO[101] = N10907 ,
      PO[102] = N10908 ,
      PO[103] = N11333 ,
      PO[104] = N11334 ,
      PO[105] = N11340 ,
      PO[106] = N11342 ,
      PO[107] = N241_O ;

   // instantiate the design into the testbench
   c7552 dut (
      .N1(N1),
      .N5(N5),
      .N9(N9),
      .N12(N12),
      .N15(N15),
      .N18(N18),
      .N23(N23),
      .N26(N26),
      .N29(N29),
      .N32(N32),
      .N35(N35),
      .N38(N38),
      .N41(N41),
      .N44(N44),
      .N47(N47),
      .N50(N50),
      .N53(N53),
      .N54(N54),
      .N55(N55),
      .N56(N56),
      .N57(N57),
      .N58(N58),
      .N59(N59),
      .N60(N60),
      .N61(N61),
      .N62(N62),
      .N63(N63),
      .N64(N64),
      .N65(N65),
      .N66(N66),
      .N69(N69),
      .N70(N70),
      .N73(N73),
      .N74(N74),
      .N75(N75),
      .N76(N76),
      .N77(N77),
      .N78(N78),
      .N79(N79),
      .N80(N80),
      .N81(N81),
      .N82(N82),
      .N83(N83),
      .N84(N84),
      .N85(N85),
      .N86(N86),
      .N87(N87),
      .N88(N88),
      .N89(N89),
      .N94(N94),
      .N97(N97),
      .N100(N100),
      .N103(N103),
      .N106(N106),
      .N109(N109),
      .N110(N110),
      .N111(N111),
      .N112(N112),
      .N113(N113),
      .N114(N114),
      .N115(N115),
      .N118(N118),
      .N121(N121),
      .N124(N124),
      .N127(N127),
      .N130(N130),
      .N133(N133),
      .N134(N134),
      .N135(N135),
      .N138(N138),
      .N141(N141),
      .N144(N144),
      .N147(N147),
      .N150(N150),
      .N151(N151),
      .N152(N152),
      .N153(N153),
      .N154(N154),
      .N155(N155),
      .N156(N156),
      .N157(N157),
      .N158(N158),
      .N159(N159),
      .N160(N160),
      .N161(N161),
      .N162(N162),
      .N163(N163),
      .N164(N164),
      .N165(N165),
      .N166(N166),
      .N167(N167),
      .N168(N168),
      .N169(N169),
      .N170(N170),
      .N171(N171),
      .N172(N172),
      .N173(N173),
      .N174(N174),
      .N175(N175),
      .N176(N176),
      .N177(N177),
      .N178(N178),
      .N179(N179),
      .N180(N180),
      .N181(N181),
      .N182(N182),
      .N183(N183),
      .N184(N184),
      .N185(N185),
      .N186(N186),
      .N187(N187),
      .N188(N188),
      .N189(N189),
      .N190(N190),
      .N191(N191),
      .N192(N192),
      .N193(N193),
      .N194(N194),
      .N195(N195),
      .N196(N196),
      .N197(N197),
      .N198(N198),
      .N199(N199),
      .N200(N200),
      .N201(N201),
      .N202(N202),
      .N203(N203),
      .N204(N204),
      .N205(N205),
      .N206(N206),
      .N207(N207),
      .N208(N208),
      .N209(N209),
      .N210(N210),
      .N211(N211),
      .N212(N212),
      .N213(N213),
      .N214(N214),
      .N215(N215),
      .N216(N216),
      .N217(N217),
      .N218(N218),
      .N219(N219),
      .N220(N220),
      .N221(N221),
      .N222(N222),
      .N223(N223),
      .N224(N224),
      .N225(N225),
      .N226(N226),
      .N227(N227),
      .N228(N228),
      .N229(N229),
      .N230(N230),
      .N231(N231),
      .N232(N232),
      .N233(N233),
      .N234(N234),
      .N235(N235),
      .N236(N236),
      .N237(N237),
      .N238(N238),
      .N239(N239),
      .N240(N240),
      .N242(N242),
      .N245(N245),
      .N248(N248),
      .N251(N251),
      .N254(N254),
      .N257(N257),
      .N260(N260),
      .N263(N263),
      .N267(N267),
      .N271(N271),
      .N274(N274),
      .N277(N277),
      .N280(N280),
      .N283(N283),
      .N286(N286),
      .N289(N289),
      .N293(N293),
      .N296(N296),
      .N299(N299),
      .N303(N303),
      .N307(N307),
      .N310(N310),
      .N313(N313),
      .N316(N316),
      .N319(N319),
      .N322(N322),
      .N325(N325),
      .N328(N328),
      .N331(N331),
      .N334(N334),
      .N337(N337),
      .N340(N340),
      .N343(N343),
      .N346(N346),
      .N349(N349),
      .N352(N352),
      .N355(N355),
      .N358(N358),
      .N361(N361),
      .N364(N364),
      .N367(N367),
      .N382(N382),
      .N241_I(N241_I),
      .N387(N387),
      .N388(N388),
      .N478(N478),
      .N482(N482),
      .N484(N484),
      .N486(N486),
      .N489(N489),
      .N492(N492),
      .N501(N501),
      .N505(N505),
      .N507(N507),
      .N509(N509),
      .N511(N511),
      .N513(N513),
      .N515(N515),
      .N517(N517),
      .N519(N519),
      .N535(N535),
      .N537(N537),
      .N539(N539),
      .N541(N541),
      .N543(N543),
      .N545(N545),
      .N547(N547),
      .N549(N549),
      .N551(N551),
      .N553(N553),
      .N556(N556),
      .N559(N559),
      .N561(N561),
      .N563(N563),
      .N565(N565),
      .N567(N567),
      .N569(N569),
      .N571(N571),
      .N573(N573),
      .N582(N582),
      .N643(N643),
      .N707(N707),
      .N813(N813),
      .N881(N881),
      .N882(N882),
      .N883(N883),
      .N884(N884),
      .N885(N885),
      .N889(N889),
      .N945(N945),
      .N1110(N1110),
      .N1111(N1111),
      .N1112(N1112),
      .N1113(N1113),
      .N1114(N1114),
      .N1489(N1489),
      .N1490(N1490),
      .N1781(N1781),
      .N10025(N10025),
      .N10101(N10101),
      .N10102(N10102),
      .N10103(N10103),
      .N10104(N10104),
      .N10109(N10109),
      .N10110(N10110),
      .N10111(N10111),
      .N10112(N10112),
      .N10350(N10350),
      .N10351(N10351),
      .N10352(N10352),
      .N10353(N10353),
      .N10574(N10574),
      .N10575(N10575),
      .N10576(N10576),
      .N10628(N10628),
      .N10632(N10632),
      .N10641(N10641),
      .N10704(N10704),
      .N10706(N10706),
      .N10711(N10711),
      .N10712(N10712),
      .N10713(N10713),
      .N10714(N10714),
      .N10715(N10715),
      .N10716(N10716),
      .N10717(N10717),
      .N10718(N10718),
      .N10729(N10729),
      .N10759(N10759),
      .N10760(N10760),
      .N10761(N10761),
      .N10762(N10762),
      .N10763(N10763),
      .N10827(N10827),
      .N10837(N10837),
      .N10838(N10838),
      .N10839(N10839),
      .N10840(N10840),
      .N10868(N10868),
      .N10869(N10869),
      .N10870(N10870),
      .N10871(N10871),
      .N10905(N10905),
      .N10906(N10906),
      .N10907(N10907),
      .N10908(N10908),
      .N11333(N11333),
      .N11334(N11334),
      .N11340(N11340),
      .N11342(N11342),
      .N241_O(N241_O)   );


   integer errshown;
   event measurePO;
   always @ measurePO begin
      if (((XPCT&MASK) !== (ALLPOS&MASK)) || (XPCT !== (~(~XPCT)))) begin
         errshown = 0;
         for (bit = 0; bit < NOUTPUTS; bit=bit + 1) begin
            if (MASK[bit]==1'b1) begin
               if (XPCT[bit] !== ALLPOS[bit]) begin
                  if (errshown==0) $display("\n// *** ERROR during capture pattern %0d, T=%t", pattern, $time);
                  $display("  %0d %0s (exp=%b, got=%b)", pattern, POnames[bit], XPCT[bit], ALLPOS[bit]);
                  nofails = nofails + 1; errshown = 1;
               end
            end
         end
      end
   end

   event forcePI_default_WFT;
   always @ forcePI_default_WFT begin
      PI = ALLPIS;
   end
   event measurePO_default_WFT;
   always @ measurePO_default_WFT begin
      #40;
      ALLPOS = PO;
      #0; #0 -> measurePO;
      `ifdef tmax_iddq
         #0; ->IDDQ;
      `endif
   end

   always @ IDDQ begin
   `ifdef tmax_iddq
      $ssi_iddq("strobe_try");
      $ssi_iddq("status drivers leaky AAA_tmax_testbench_1_16.leaky");
   `endif
   end

   event capture;
   always @ capture begin
      ->forcePI_default_WFT;
      #100; ->measurePO_default_WFT;
   end


   initial begin

      //
      // --- establish a default time format for %t
      //
      $timeformat(-9,2," ns",18);

      //
      // --- default verbosity to 2 but also allow user override by
      //     using '+define+tmax_msg=N' on verilog compile line.
      //
      `ifdef tmax_msg
         verbose = `tmax_msg ;
      `else
         verbose = 2 ;
      `endif

      //
      // --- default pattern reporting interval to 5 but also allow user
      //     override by using '+define+tmax_rpt=N' on verilog compile line.
      //
      `ifdef tmax_rpt
         report_interval = `tmax_rpt ;
      `else
         report_interval = 5 ;
      `endif

      //
      // --- support generating Extened VCD output by using
      //     '+define+tmax_vcde' on verilog compile line.
      //
      `ifdef tmax_vcde
         // extended VCD, see IEEE Verilog P1364.1-1999 Draft 2
         if (verbose >= 2) $display("// %t : opening Extended VCD output file", $time);
         $dumpports( dut, "sim_vcde.out");
      `endif

      //
      // --- IDDQ PLI initialization
      //     User may activite by using '+define+tmax_iddq' on verilog compile line.
      //     Or by defining `tmax_iddq in this file.
      //
      `ifdef tmax_iddq
         if (verbose >= 3) $display("// %t : Initializing IDDQ PLI", $time);
         $ssi_iddq("dut AAA_tmax_testbench_1_16.dut");
         $ssi_iddq("verb on");
         $ssi_iddq("cycle 0");
         //
         // --- User may select one of the following two methods for fault seeding:
         //     #1 faults seeded by PLI (default)
         //     #2 faults supplied in a file
         //     Comment out the unused lines as needed (precede with '//').
         //     Replace the 'FAULTLIST_FILE' string with the actual file pathname.
         //
         $ssi_iddq("seed SA AAA_tmax_testbench_1_16.dut");   // no file, faults seeded by PLI
         //
         // $ssi_iddq("scope AAA_tmax_testbench_1_16.dut");   // set scope for faults from a file
         // $ssi_iddq("read_tmax FAULTLIST_FILE"); // read faults from a file
         //
      `endif

      POnames[0] = "N387";
      POnames[1] = "N388";
      POnames[2] = "N478";
      POnames[3] = "N482";
      POnames[4] = "N484";
      POnames[5] = "N486";
      POnames[6] = "N489";
      POnames[7] = "N492";
      POnames[8] = "N501";
      POnames[9] = "N505";
      POnames[10] = "N507";
      POnames[11] = "N509";
      POnames[12] = "N511";
      POnames[13] = "N513";
      POnames[14] = "N515";
      POnames[15] = "N517";
      POnames[16] = "N519";
      POnames[17] = "N535";
      POnames[18] = "N537";
      POnames[19] = "N539";
      POnames[20] = "N541";
      POnames[21] = "N543";
      POnames[22] = "N545";
      POnames[23] = "N547";
      POnames[24] = "N549";
      POnames[25] = "N551";
      POnames[26] = "N553";
      POnames[27] = "N556";
      POnames[28] = "N559";
      POnames[29] = "N561";
      POnames[30] = "N563";
      POnames[31] = "N565";
      POnames[32] = "N567";
      POnames[33] = "N569";
      POnames[34] = "N571";
      POnames[35] = "N573";
      POnames[36] = "N582";
      POnames[37] = "N643";
      POnames[38] = "N707";
      POnames[39] = "N813";
      POnames[40] = "N881";
      POnames[41] = "N882";
      POnames[42] = "N883";
      POnames[43] = "N884";
      POnames[44] = "N885";
      POnames[45] = "N889";
      POnames[46] = "N945";
      POnames[47] = "N1110";
      POnames[48] = "N1111";
      POnames[49] = "N1112";
      POnames[50] = "N1113";
      POnames[51] = "N1114";
      POnames[52] = "N1489";
      POnames[53] = "N1490";
      POnames[54] = "N1781";
      POnames[55] = "N10025";
      POnames[56] = "N10101";
      POnames[57] = "N10102";
      POnames[58] = "N10103";
      POnames[59] = "N10104";
      POnames[60] = "N10109";
      POnames[61] = "N10110";
      POnames[62] = "N10111";
      POnames[63] = "N10112";
      POnames[64] = "N10350";
      POnames[65] = "N10351";
      POnames[66] = "N10352";
      POnames[67] = "N10353";
      POnames[68] = "N10574";
      POnames[69] = "N10575";
      POnames[70] = "N10576";
      POnames[71] = "N10628";
      POnames[72] = "N10632";
      POnames[73] = "N10641";
      POnames[74] = "N10704";
      POnames[75] = "N10706";
      POnames[76] = "N10711";
      POnames[77] = "N10712";
      POnames[78] = "N10713";
      POnames[79] = "N10714";
      POnames[80] = "N10715";
      POnames[81] = "N10716";
      POnames[82] = "N10717";
      POnames[83] = "N10718";
      POnames[84] = "N10729";
      POnames[85] = "N10759";
      POnames[86] = "N10760";
      POnames[87] = "N10761";
      POnames[88] = "N10762";
      POnames[89] = "N10763";
      POnames[90] = "N10827";
      POnames[91] = "N10837";
      POnames[92] = "N10838";
      POnames[93] = "N10839";
      POnames[94] = "N10840";
      POnames[95] = "N10868";
      POnames[96] = "N10869";
      POnames[97] = "N10870";
      POnames[98] = "N10871";
      POnames[99] = "N10905";
      POnames[100] = "N10906";
      POnames[101] = "N10907";
      POnames[102] = "N10908";
      POnames[103] = "N11333";
      POnames[104] = "N11334";
      POnames[105] = "N11340";
      POnames[106] = "N11342";
      POnames[107] = "N241_O";
      nofails = 0; pattern = -1; lastpattern = 0;
      prev_pat = -2; error_banner = -2;
      /*** No test setup procedure ***/


      /*** Non-scan test ***/

      if (verbose >= 1) $display("// %t : Begin patterns, first pattern = 0", $time);
pattern = 0; // 0
ALLPIS = 207'b110100001001000011010010110100000010110110011110000101111111110010111111100101111101000101110111010010101100110000001000010010101010001110110010011011000011101010100110011110001100001101001000001011100110101;
XPCT = 108'b111011110110000110100100000111100110100011111111111111011111110010011111010111000001110011111111001100111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 200

pattern = 1; // 200
ALLPIS = 207'b111010000100100001101001011010000001011011001111000010111111111001011111110010111110100010111011101001010110011000000100001001010101000111011001001101100001110101010011001111000110000110100100000101110011010;
XPCT = 108'b111001110011000011010010000001110011010111111101011011000000111100001010000010010111100111000110110010101110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 400

pattern = 2; // 400
ALLPIS = 207'b101001001011010011100110011001000010011011111001100100100000001110010000011100100010010100101010100110000111111100001010010110000000101101011110111101110011010000001111111001101111001110011010001001011111000;
XPCT = 108'b111111001111100111001101000101011111110001101100101111011111100110111111010100110111110101111000011110010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 600

pattern = 3; // 600
ALLPIS = 207'b000000101100101010100001111000100011111011100010110111101111110101110111101011101100001111100010000001101111001110001101011001101010011000011101000101111010000010100001100010111011101010000101001111001001001;
XPCT = 108'b000100011101110101000010100111001001111101111011110100001111010110110101101111011100111001000000111100111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 800

pattern = 4; // 800
ALLPIS = 207'b010100011111010110000010001000010011001011101111011110001000001000000100010000001011000010000110010010011011010111001110111110011111000010111100111001111110101011110110101111010001111000001010101100000010001;
XPCT = 108'b001101110000111100000101010100000010101110111001111110011111011000111111110100000110111000111110110001110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1000

pattern = 5; // 1000
ALLPIS = 207'b001010001111101011000001000100001001100101110111101111000100000100000010001000000101100001000011001001001101101011100111011111001111100001011110011100111111010101111011010111101000111100000101010110000001000;
XPCT = 108'b001010111100011110000010101010000001010101111010001010001111000100101111100101101001110000111110111101101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1200

pattern = 6; // 1200
ALLPIS = 207'b110001001110110110110010010110000110000100100101110010011101110000111110100001111111110101010110110110001010000101111011111101001101111110011101010101011100000000011011110101111000010011001010100000100110001;
XPCT = 108'b111110101100001001100101010000100110111011111101111111011111101110101111001111010100110101000000001111100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1400

pattern = 7; // 1400
ALLPIS = 207'b111000100111011011011001001011000011000010010010111001001110111000011111010000111111111010101011011011000101000010111101111110100110111111001110101010101110000000001101111010111100001001100101010000010011000;
XPCT = 108'b110111011110000100110010101000010011111011111111111111101111101001011111000110110000111011011110111111111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1600

pattern = 8; // 1600
ALLPIS = 207'b001000011010101110111110010001100011010111010111011001011000101110110000001101100010111000100010111111001110010001010110101101111001010001010101001110010100101010100000100011010010001001111010100011101111001;
XPCT = 108'b000100010001000100111101010011101111101011011011110100011111101100001111011100111100111011000001000111000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1800

pattern = 9; // 1800
ALLPIS = 207'b000100001101010111011111001000110001101011101011101100101100010111011000000110110001011100010001011111100111001000101011010110111100101000101010100111001010010101010000010001101001000100111101010001110111100;
XPCT = 108'b000010001100100010011110101001110111100011111001111110001111001001001111110100101011110111111110011011101110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2000

pattern = 10; // 2000
ALLPIS = 207'b100010000110101011101111100100011000110101110101110110010110001011101100000011011000101110001000101111110011100100010101101011011110010100010101010011100101001010101000001000110100100010011110101000111011110;
XPCT = 108'b110001001010010001001111010100111011001011111100001011111001101001010100010110100111111110000000010011001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2200

pattern = 11; // 2200
ALLPIS = 207'b000101001010010110100101000110001110101100100100111110110100110111001001100100010001010010110011000101010101000010000010100111000101000100111000110010110001001111110010011010010110011100000111011111111011010;
XPCT = 108'b001011010011001110000011101111111011101101111001111110010000011010011110010010100110100010100110010010101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2400

pattern = 12; // 2400
ALLPIS = 207'b010110101100001000000000010111000101100000001100011010100101101001011011010111110101101100101110110000000110010001001001000001001000101100101110000010011011001101011111010011000111000011001011100100011011000;
XPCT = 108'b001010010011100001100101110000011011010111111001011010001111100010101111101111111011111110000000110110110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2600

pattern = 13; // 2600
ALLPIS = 207'b001011010110000100000000001011100010110000000110001101010010110100101101101011111010110110010111011000000011001000100100100000100100010110010111000001001101100110101111101001100011100001100101110010001101100;
XPCT = 108'b001101001001110000110010111010001101010001111010001010000000110101111110110011101101101101111111111000001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2800

pattern = 14; // 2800
ALLPIS = 207'b010001100010000001010010110001110011101110011101000011010110101000101001010000000000011110111100111110101101010100011010000010111000000101111001111011100101011001110001101010111101111101111010110010100000011;
XPCT = 108'b000101011110111110111101011010100000111011111011111110010000000110001110101001001011100000000110110011111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3000

pattern = 15; // 3000
ALLPIS = 207'b001000110001000000101001011000111001110111001110100001101011010100010100101000000000001111011110011111010110101010001101000001011100000010111100111101110010101100111000110101011110111110111101011001010000001;
XPCT = 108'b000110100111011111011110101101010000101011111010101110011111011010010101110100011000110000011110110111111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3200

pattern = 16; // 3200
ALLPIS = 207'b110000010001100011000110011000011110001101111001010101001010011000110101110001111101000010011000011101000111100101001110110010000100001111101100000101111010111100111010000100100011010010010110100111001110101;
XPCT = 108'b111000101001101001001011010011001110100110111111111111011111100000101111010111111101111100011110011100111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3400

pattern = 17; // 3400
ALLPIS = 207'b101100000001110010110001111000001101110000100010101111011010111110100101011101000011100100111011011100001111000010101111001011101000001001000100011001111110110100111011011100011101100100000011011000000001111;
XPCT = 108'b111011100110110010000001101100000001111000111110101111011001100000111110000101110001110110100110101100001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3600

pattern = 18; // 3600
ALLPIS = 207'b110110000000111001011000111100000110111000010001010111101101011111010010101110100001110010011101101110000111100001010111100101110100000100100010001100111111011010011101101110001110110010000001101100000000111;
XPCT = 108'b110101110111011001000000110100000000010111111111011011010000100010011110100000010100101100000111110000011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3800

pattern = 19; // 3800
ALLPIS = 207'b111011000000011100101100011110000011011100001000101011110110101111101001010111010000111001001110110111000011110000101011110010111010000010010001000110011111101101001110110111000111011001000000110110000000011;
XPCT = 108'b111110110011101100100000011010000000000111111111011011110110110000101111001000100010100110100110100010001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4000

pattern = 20; // 4000
ALLPIS = 207'b011101100000001110010110001111000001101110000100010101111011010111110100101011101000011100100111011011100001111000010101111001011101000001001000100011001111110110100111011011100011101100100000011011000000001;
XPCT = 108'b001011011001110110010000001111000000110011111011111110010000010001111110101001000001100010111110000001000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4200

pattern = 21; // 4200
ALLPIS = 207'b101110110000000111001011000111100000110111000010001010111101101011111010010101110100001110010011101101110000111100001010111100101110100000100100010001100111111011010011101101110001110110010000001101100000000;
XPCT = 108'b111101101000111011001000000101100000011111111101010001110000101100111110100010110110100100111111110101101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4400

pattern = 22; // 4400
ALLPIS = 207'b100011010001000000110111010111110010101101111111000000100001000111000010101111000111000010111110100100010100101110001101001100111101011110100000010011110000010111001111101000110100110110000000001101010110101;
XPCT = 108'b111101001010011011000000000101010110011101111100001011001111011100011111111101000000110001111111000101000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4600

pattern = 23; // 4600
ALLPIS = 207'b000101100001100011001001011111111011100000100001100101101111010001011110110010011110100100101000000000100110100111001110110100110100100001100010010010111011100001000001101010010110010110001000001101001101111;
XPCT = 108'b000101010011001011000100000101001101111111111011111110001001110111011110011101111010111111100001111110100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4800

pattern = 24; // 4800
ALLPIS = 207'b110110111001110010110110011011111111000110001110110111001000011010010000111100110010010111100011010010111111100011101111001000110000011110000011010010011110011010000110101011000111000110001100001101000000010;
XPCT = 108'b111101010011100011000110000101000000000111111111011011001111001110101111111110100100110110000110100100000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5000

pattern = 25; // 5000
ALLPIS = 207'b011011011100111001011011001101111111100011000111011011100100001101001000011110011001001011110001101001011111110001110111100100011000001111000001101001001111001101000011010101100011100011000110000110100000001;
XPCT = 108'b001010101001110001100011000010100000010111101011011010011111010010111111111111010101110111100000011011000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5200

pattern = 26; // 5200
ALLPIS = 207'b011001100111011111111111010010111101000111111101101000001101110100011011101010110001100000001111100110000011001000110011100000100110001001010010101111100100001100000111110100111101111100101011001000110110101;
XPCT = 108'b001110101110111110010101100100110110111011111001111110001111011111011111000101101111111011111000010010000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5400

pattern = 27; // 5400
ALLPIS = 207'b101100110011101111111111101001011110100011111110110100000110111010001101110101011000110000000111110011000001100100011001110000010011000100101001010111110010000110000011111010011110111110010101100100011011010;
XPCT = 108'b111111010111011111001010110000011011111111111101111111001001110000111110001100000010110001000000110000000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5600

pattern = 28; // 5600
ALLPIS = 207'b000010010000110100101101000000101101100111100001011111111100101111111001011111010001011101110100101011001100000010000100101010100011101100100110110000111010101001100111100011000011010010000010111001101011000;
XPCT = 108'b001100010001101001000001011101101011010011111011010000001111101000101111100100011100111101000000001011101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5800

pattern = 29; // 5800
ALLPIS = 207'b100001001000011010010110100000010110110011110000101111111110010111111100101111101000101110111010010101100110000001000010010101010001110110010011011000011101010100110011110001100001101001000001011100110101100;
XPCT = 108'b111110001000110100100000101100110101110101111111110101101001010010111110100100000010111001000001011001000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6000

pattern = 30; // 6000
ALLPIS = 207'b010000100100001101001011010000001011011001111000010111111111001011111110010111110100010111011101001010110011000000100001001010101000111011001001101100001110101010011001111000110000110100100000101110011010110;
XPCT = 108'b000111001000011010010000010110011010111111111011111110001001101101111110101111000000110100100000100000111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6200

pattern = 31; // 6200
ALLPIS = 207'b101000010010000110100101101000000101101100111100001011111111100101111111001011111010001011101110100101011001100000010000100101010100011101100100110110000111010101001100111100011000011010010000010111001101011;
XPCT = 108'b110111100100001101001000001011001101101101111110100101110000011111011110010011010000101001011111101100100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6400

pattern = 32; // 6400
ALLPIS = 207'b100011001100100001000000010011010110001010010101001001111100011010011000001111011001110100100110011111111100000000100100010100101101110111000101111000010011101110111011111110101111001110110100111111110000001;
XPCT = 108'b111111111111100111011010011111110000010101111110001011010000001000101110101010101101100000111111000011000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6600

pattern = 33; // 6600
ALLPIS = 207'b110001100110010000100000001001101011000101001010100100111110001101001100000111101100111010010011001111111110000000010010001010010110111011100010111100001001110111011101111111010111100111011010011111111000000;
XPCT = 108'b110111110011110011101101001111111000111111111101111111111001000011101110100111010001110100000001100100100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6800

pattern = 34; // 6800
ALLPIS = 207'b111011111111101001010000010111100011101000110000011011100011011100111110001100101111101001101111111000000011000000101101010001100110101010110100100110010111010101010101000001000100111101011001110000001100001;
XPCT = 108'b110000000010011110101100111000001100010011111111011011111111111011100111010111011000110011111110101111101001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7000

pattern = 35; // 7000
ALLPIS = 207'b111110110011010101101000011000100111111110001101000100001101110100000111001001001110000000010001100011111101100000110010111100011110100010011111101011011000000100010001011110001101010000011000000111110110001;
XPCT = 108'b110011110110101000001100000011110110010111111101011011011111111110111111100101110011111101011000001111000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7200

pattern = 36; // 7200
ALLPIS = 207'b101110001010100101111010001111100010111010101001110101111101010000001101110101111111011010010111010111000001011000011110100101010001010011000101000110111111110110011001101000110100110011011100011110000101100;
XPCT = 108'b110101001010011001101110001110000101011110011110001011100000001111111110000001010100101101111110000001100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7400

pattern = 37; // 7400
ALLPIS = 207'b110100001001110011111101010100100111010111000001110011000010110010011110110101100110011001101101110100011100101100101011000110000101011110100111011011001100010101110111001010110101010111011010110000110010111;
XPCT = 108'b111001011010101011101101011000110010111011011111111111101111001101010101100100100101110101000110110101110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7600

pattern = 38; // 7600
ALLPIS = 207'b111110001110111101111111000110011111111111100101010101001100110110111111100010000000010010111101000010111011001011101110100101001100100000101100001110100000101011100110001100000010011011000010010011111100100;
XPCT = 108'b111001100001001101100001001011111100000011111111011011000000000101011110110000110101101010111111011001100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7800

pattern = 39; // 7800
ALLPIS = 207'b111111000111011110111111100011001111111111110010101010100110011011011111110001000000001001011110100001011101100101110111010010100110010000010110000111010000010101110011000110000001001101100001001001111110010;
XPCT = 108'b111000110000100110110000100101111110010010111101011011110000001111111110000010001111100011111111000000001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8000

pattern = 40; // 8000
ALLPIS = 207'b011111100011101111011111110001100111111111111001010101010011001101101111111000100000000100101111010000101110110010111011101001010011001000001011000011101000001010111001100011000000100110110000100100111111001;
XPCT = 108'b000100010000010011011000010000111111010111101011011010011111011011001111000100001100110111111000110110000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8200

pattern = 41; // 8200
ALLPIS = 207'b101100111101010110101111101011100101110101101001100011010101111100101111110011001001110110110001110111101011011001111001100000000100010011000000011001100111101011100111001111001111011101101100101101101111101;
XPCT = 108'b111001110111101110110110010101101111110111111111111111011111000100001111001110000101110001011001110111010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8400

pattern = 42; // 8400
ALLPIS = 207'b110101010010001010010111100110100100110000100001111000010110100100001111110110111101001111111110100100001001101100011000100100101111111110100101110100100000011011001000011001001000100000000010101001000111111;
XPCT = 108'b110011000100010000000001010101000111100011111101111111100000101111001110110010111110101010111110001100111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8600

pattern = 43; // 8600
ALLPIS = 207'b011010101001000101001011110011010010011000010000111100001011010010000111111011011110100111111111010010000100110110001100010010010111111111010010111010010000001101100100001100100100010000000001010100100011111;
XPCT = 108'b000001101010001000000000101000100011000111111001011010001111010100001111011110010111111101011001111111100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8800

pattern = 44; // 8800
ALLPIS = 207'b101110011000000011100101101010111111000110011101010111111001110011011011110010110110100111011001110110111110011011100010011101100110001000101100100101011011101000001001111000111101000110110100010101100001110;
XPCT = 108'b110111001110100011011010001001100001011101111110001011000000000000111010100010100000100111011111100011111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9000

pattern = 45; // 9000
ALLPIS = 207'b110111001100000001110010110101011111100011001110101011111100111001101101111001011011010011101100111011011111001101110001001110110011000100010110010010101101110100000100111100011110100011011010001010110000111;
XPCT = 108'b110111100111010001101101000110110000001011111111011011000000111001011110001001000010100100011000101100011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9200

pattern = 46; // 9200
ALLPIS = 207'b001111011001110001111100110111101010110111101100000111111101011001001111010110100011111010001110011110110101110011101010001101010111111101100010100000110001000100100111001110111111000001011000000010100100000;
XPCT = 108'b001001111111100000101100000010100100011011111011011010011111110100110111101100110101111111011001011011100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9400

pattern = 47; // 9400
ALLPIS = 207'b100111101100111000111110011011110101011011110110000011111110101100100111101011010001111101000111001111011010111001110101000110101011111110110001010000011000100010010011100111011111100000101100000001010010000;
XPCT = 108'b111100110111110000010110000001010010011011111111011011111111010000011111001100101000111011000000110000010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9600

pattern = 48; // 9600
ALLPIS = 207'b110011110110011100011111001101111010101101111011000001111111010110010011110101101000111110100011100111101101011100111010100011010101111111011000101000001100010001001001110011101111110000010110000000101001000;
XPCT = 108'b110110011111111000001011000000101001010011111111011011111001011011111010100110000110110010000000100100101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9800

pattern = 49; // 9800
ALLPIS = 207'b111001111011001110001111100110111101010110111101100000111111101011001001111010110100011111010001110011110110101110011101010001101010111111101100010100000110001000100100111001110111111000001011000000010100100;
XPCT = 108'b110111001011111100000101100000010100101011111101111111101111010001011111111101010001110011111111100111001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10000

pattern = 50; // 10000
ALLPIS = 207'b111101010010010010100011101010111001011111111010010001110011100000101010010001110100110011010010000011000001101011000011000000110111011000111110111101010010001100110010110000110010110000110110001111110101000;
XPCT = 108'b111110001001011000011011000111110101101110111111111111010000000001111110111011111000101100011111110000001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10200

pattern = 51; // 10200
ALLPIS = 207'b001101111110010101001000100000010011011000100001001001011110101111011110101100101000000010000001110000110010011010000110101110110110111010101000101011001110111010101010101101110100000101100011000011110101011;
XPCT = 108'b001101101010000010110001100011110101101011111010101110010000100010000110110011010100100111111001100011100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10400

pattern = 52; // 10400
ALLPIS = 207'b000110111111001010100100010000001001101100010000100100101111010111101111010110010100000001000000111000011001001101000011010111011011011101010100010101100111011101010101010110111010000010110001100001111010101;
XPCT = 108'b000010111101000001011000110001111010011001011001011010001111010010011111000110011011111111111111010110110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10600

pattern = 53; // 10600
ALLPIS = 207'b000000010011000100010010011011010010111100011101011011101011110001101111100100010011110100000110000011110000100110000101111111000000011001101111110010100000000000010001010101110010001111101100001111001101011;
XPCT = 108'b000010101001000111110110000111001101111101111011111110001111110000001111001110111001110011011000000001000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10800

pattern = 54; // 10800
ALLPIS = 207'b110011001000010000000100110101100010100101010010011111000110100110000011110110011101001001100111111111000000001001000101001011011101110001011110000100111011101110111111101011110011101101001111111100000011011;
XPCT = 108'b111101011001110110100111111100000011011111111111011011110110000111111111010000001001101100100110011110011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11000

pattern = 55; // 11000
ALLPIS = 207'b011001100100001000000010011010110001010010101001001111100011010011000001111011001110100100110011111111100000000100100010100101101110111000101111000010011101110111011111110101111001110110100111111110000001101;
XPCT = 108'b001110101100111011010011111110000001111111111011111110000000111001111110000001011011100001111110000010000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11200

pattern = 56; // 11200
ALLPIS = 207'b001100110010000100000001001101011000101001010100100111110001101001100000111101100111010010011001111111110000000010010001010010110111011100010111100001001110111011101111111010111100111011010011111111000000110;
XPCT = 108'b001111011110011101101001111111000000111101011010101110010000101110100100001011010000101000000110000110110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11400

pattern = 57; // 11400
ALLPIS = 207'b000110011001000010000000100110101100010100101010010011111000110100110000011110110011101001001100111111111000000001001000101001011011101110001011110000100111011101110111111101011110011101101001111111100000011;
XPCT = 108'b001111100111001110110100111111100000011101111011010000001111010101101111000100000000110001111001010111100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11600

pattern = 58; // 11600
ALLPIS = 207'b101101101111010111111110010100111110111110000001000010000010001001100010000110001011000111100110011001100101101100100000000000011011101011111011011101001000011111000110001110011100010101101110100001111010110;
XPCT = 108'b111001110110001010110111010001111010101011111101111111000110001011001111110011110111100101011111111011101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11800

pattern = 59; // 11800
ALLPIS = 207'b110110110111101011111111001010011111011111000000100001000001000100110001000011000101100011110011001100110010110110010000000000001101110101111101101110100100001111100011000111001110001010110111010000111101011;
XPCT = 108'b111000110111000101011011101000111101010011111111011011001111101110001111100100101101111011100001011011100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12000

pattern = 60; // 12000
ALLPIS = 207'b100011011010111010010000100001011110111010101100111011110101110011110110110110011010011100111001010101010100001011100101000000001000100101001011110100100101011011010100011001000110010101101010010001101111010;
XPCT = 108'b110011000011001010110101001001101111000001111111010001110000010111001110100000110110101111011111110111101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12200

pattern = 61; // 12200
ALLPIS = 207'b010010101111110101010011110101111010100110110100110101111100000101100100010001011010100101111000110101010110010110110100101000011100010101101100110100111110110011101101001110110011100010011000011011101001100;
XPCT = 108'b000001111001110001001100001111101001011011111011011010011111111101001111101111000101111101011111011010111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12400

pattern = 62; // 12400
ALLPIS = 207'b001001010111111010101001111010111101010011011010011010111110000010110010001000101101010010111100011010101011001011011010010100001110001010110110011010011111011001110110100111011001110001001100001101110100110;
XPCT = 108'b001100110100111000100110000101110100101111111001110100001111110111001111011101001001111111100001011011000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12600

pattern = 63; // 12600
ALLPIS = 207'b001111111010101001010100001010010001101010110111100100101101101001001110100100000000010011001001011111001111011110010110100101011000001001010110111011101111101001011011100111101010001001111101100010100111111;
XPCT = 108'b001100111101000100111110110010100111010001111000001010000000101001111110100010101110101011000000110110110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12800

pattern = 64; // 12800
ALLPIS = 207'b011111001011110111001011010000100011011100110111101110000111000110110011010011001001110100000110110100000101001100011010110100110110010000001111011101000111100101111100110001000110000001111010100101110000100;
XPCT = 108'b000110000011000000111101010001110000000111111001011010001111111010001111011110111010111111011001111110001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13000

pattern = 65; // 13000
ALLPIS = 207'b001111100101111011100101101000010001101110011011110111000011100011011001101001100100111010000011011010000010100110001101011010011011001000000111101110100011110010111110011000100011000000111101010010111000010;
XPCT = 108'b001011001001100000011110101010111000000001110010001010011111001001001111111110000001111111011000001110110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13200

pattern = 66; // 13200
ALLPIS = 207'b001010011101101010001100100000110110001001001100111001100011111000001110110010111001011010100111110100100100111111100110101101010110001111111000101010011001100110011001000010001101110101110000001000100110111;
XPCT = 108'b000000010110111010111000000100100110010011110010001010001111000000000101000100101101110100100111011110011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13400

pattern = 67; // 13400
ALLPIS = 207'b010100010000110001011100000010010010111101010011101111011001111010110010101111101011110101011010110001111011111001101001101011011000010110000011100100000010010110000101010111101101010111101011010010110100110;
XPCT = 108'b000010111110101011110101101010110100110011111011111110000110010111111111000011011001100100000111000110110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13600

pattern = 68; // 13600
ALLPIS = 207'b001010001000011000101110000001001001011110101001110111101100111101011001010111110101111010101101011000111101111100110100110101101100001011000001110010000001001011000010101011110110101011110101101001011010011;
XPCT = 108'b001101011011010101111010110101011010001011111011011010000000110101101110110001110100101010111000100001110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13800

pattern = 69; // 13800
ALLPIS = 207'b000101000100001100010111000000100100101111010100111011110110011110101100101011111010111101010110101100011110111110011010011010110110000101100000111001000000100101100001010101111011010101111010110100101101001;
XPCT = 108'b000010101101101010111101011000101101111101101011111110010110110101001111110011001111100100011110100100010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14000

pattern = 70; // 14000
ALLPIS = 207'b000010100010000110001011100000010010010111101010011101111011001111010110010101111101011110101011010110001111011111001101001101011011000010110000011100100000010010110000101010111101101010111101011010010110100;
XPCT = 108'b000101011110110101011110101110010110001011110011011010001111010101000101010111010100111001000001110111001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14200

pattern = 71; // 14200
ALLPIS = 207'b111011110000011101100011100110100101000100111011000100011101111110100110100000010001110011111111100000110100101101000011010011000000101110101010110100100100010100001001000011111101000101110110100111100010000;
XPCT = 108'b110000011110100010111011010011100010011111111101011011011111100010111111110101011001111000100001100011010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14400

pattern = 72; // 14400
ALLPIS = 207'b011001101010100001101101101101000101111001000110001010000001000100001110010011101011111000000000000011111010010010000000011010000101010100110000111100111110111010010110100101100100111000011011111101011000001;
XPCT = 108'b001100101010011100001101111101011000100111111001111110011001001111001110001110010010110111000000001001000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14600

pattern = 73; // 14600
ALLPIS = 207'b101100110101010000110110110110100010111100100011000101000000100010000111001001110101111100000000000001111101001001000000001101000010101010011000011110011111011101001011010010110010011100001101111110101100000;
XPCT = 108'b111010011001001110000110111110101100111101111110101111111111100110111111000111101001110001011001010111010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14800

pattern = 74; // 14800
ALLPIS = 207'b011011110101111111100101001111101111100000010000100000100010011000100001100010110001111001100110011001011011001000000000000110111010111110110111010010000111110001100011100111000101011011101000011110101100110;
XPCT = 108'b001100110010101101110100001110101100010111111001011010001111110001101111000101111010110100100001100100111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15000

pattern = 75; // 15000
ALLPIS = 207'b101101111010111111110010100111110111110000001000010000010001001100010000110001011000111100110011001100101101100100000000000011011101011111011011101001000011111000110001110011100010101101110100001111010110011;
XPCT = 108'b110110011001010110111010000111010110110101111101111111110000110011101110000011001010100010000111110011100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15200

pattern = 76; // 15200
ALLPIS = 207'b011011011110101111111100101001111101111100000010000100000100010011000100001100010110001111001100110011001011011001000000000000110111010111110110111010010000111110001100011100111000101011011101000011110101100;
XPCT = 108'b000011101100010101101110100011110101001011111001011010001001000000011110010101010010111100000001011000011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15400

pattern = 77; // 15400
ALLPIS = 207'b001100001110010010100110111001011110110101011000010000101100000001101111111001011000110100101000000110101011000000001100101001101010100011101001100010110001100110010110011100010001101100001110100111010001100;
XPCT = 108'b001011100000110110000111010011010001101100111001111110000000010110111110011011110011100010011110110001000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15600

pattern = 78; // 15600
ALLPIS = 207'b101011110100001100101100100000000111110011101111111011100111100010001010001000001110000001001001001000011101111000010010001011000111100001010011011010011100010101000011011001011000001111110101001110100000011;
XPCT = 108'b111011000100000111111010100110100000011111111111011011010000100111101110011011010110100100011110100110110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15800

pattern = 79; // 15800
ALLPIS = 207'b110101111010000110010110010000000011111001110111111101110011110001000101000100000111000000100100100100001110111100001001000101100011110000101001101101001110001010100001101100101100000111111010100111010000001;
XPCT = 108'b110101101110000011111101010011010000110111101111111111010000001000111110010001000110101000011110010011010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16000

pattern = 80; // 16000
ALLPIS = 207'b100001010000110011000011011101011110001011000101101111110000111101111110101000011001000100100001001111101000101111001110111000110010011111100011111001100010000100111110000111011010101101110000001110100101100;
XPCT = 108'b111000110101010110111000000110100101101101111110100101001111000110001111011101001011110100100000011010111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16200

pattern = 81; // 16200
ALLPIS = 207'b101000110100111100101100011100010010101111010010010110100000011101100000100110111101001011000000101010100010010111111110001111001100001000100010111001010010001110110011111011001110001110100101001001110001110;
XPCT = 108'b111111010111000111010010100101110001110011111101111111110000010110111110001000010010100011111000000111001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16400

pattern = 82; // 16400
ALLPIS = 207'b010100011010011110010110001110001001010111101001001011010000001110110000010011011110100101100000010101010001001011111111000111100110000100010001011100101001000111011001111101100111000111010010100100111000111;
XPCT = 108'b000111101011100011101001010000111000110111111011111110010000100000011110000010100000100110111110000010011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16600

pattern = 83; // 16600
ALLPIS = 207'b001010001101001111001011000111000100101011110100100101101000000111011000001001101111010010110000001010101000100101111111100011110011000010001000101110010100100011101100111110110011100011101001010010011100011;
XPCT = 108'b000111111001110001110100101010011100001011111010001010001111101101001111111111110000111101000001111101010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16800

pattern = 84; // 16800
ALLPIS = 207'b000001110000111100001011101100011001001111100101111111010011100011101110010000101101000011000101001111000011110010001011110011110101110010010101001110101110110100001100100010010100111011010111010001110110011;
XPCT = 108'b000100010010011101101011101001110110101011111010101110010000100111111010001010100110101011111001111110100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17000

pattern = 85; // 17000
ALLPIS = 207'b110100011100110000001010010110000000010110010100011110001110011110101101111001101100110101100000100010000101011110000100100100100001001010101000001110100111011100011011000000100000010011001001010011111100010;
XPCT = 108'b111000001000001001100100101011111100110011111101111111011001011001001110000111111111111101100001000111001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17200

pattern = 86; // 17200
ALLPIS = 207'b011001100110101011011011000001110101011111111110100101101010001100101110100110010000110001001101101011011111000101001011111110011011000101110000001111011100001101100110111111110010010100000000100000100001011;
XPCT = 108'b001111111001001010000000010000100001101011110011111110010000110011001110010010110111101110100001010100011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17400

pattern = 87; // 17400
ALLPIS = 207'b001010010111111000010000001001000011100010100111111001110110100010100100010000111100111000111011011100011100110001011110010110001100010010110101100001000110100101001111110011101101001001001110101111011001110;
XPCT = 108'b001110011110100100100111010111011001010101111010001010001111011011001111000111101000111010000111111000101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17600

pattern = 88; // 17600
ALLPIS = 207'b111101010111011001000101110110011100011011100011011101100011010010001101111010101111110101001101100011011000011000110110011000010011001110001001110101000000011110001011000001010101111100111010011001001111111;
XPCT = 108'b111000000010111110011101001101001111111011111111111111001111011110001111100111001101110000011000011100001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17800

pattern = 89; // 17800
ALLPIS = 207'b111110101011101100100010111011001110001101110001101110110001101001000110111101010111111010100110110001101100001100011011001100001001100111000100111010100000001111000101100000101010111110011101001100100111111;
XPCT = 108'b110100001101011111001110100100100111010111111101011011111111111101101111001111001110110000111001000111111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18000

pattern = 90; // 18000
ALLPIS = 207'b000111001001010011011100101111011010101100001000010110000000110111111100101100011010010100000011010101100000000110010100110101010001110100110001011000110011001011001110001000110110000111010011101000110000111;
XPCT = 108'b001001001011000011101001110100110000001011111000000000001111100101011111001101001011111001011001100010001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18200

pattern = 91; // 18200
ALLPIS = 207'b000011100100101001101110010111101101010110000100001011000000011011111110010110001101001010000001101010110000000011001010011010101000111010011000101100011001100101100111000100011011000011101001110100011000011;
XPCT = 108'b001000100101100001110100111000011000011111111011010000010000111101111110101011110111100111111110011000110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18400

pattern = 92; // 18400
ALLPIS = 207'b110000111001001010011011100101111011010101100001000010110000000110111111100101100011010010100000011010101100000000110010100110101010001110100110001011000110011001011001110001000110110000111010011101000110000;
XPCT = 108'b110110000011011000011101001101000110110111111101111111011111011111011111100110011010111100011110101001001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18600

pattern = 93; // 18600
ALLPIS = 207'b011110111100111101001010001011111011111001111100011101011001010000111111110000011100000011111010001000110101111000101101000001000111011010000100101110000100010111100010001101110110111000000101100011100111100;
XPCT = 108'b001001101011011100000010110011100111001011111011011010010000111100011110010000010101101001111110100000000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18800

pattern = 94; // 18800
ALLPIS = 207'b001111011110011110100101000101111101111100111110001110101100101000011111111000001110000001111101000100011010111100010110100000100011101101000010010111000010001011110001000110111011011100000010110001110011110;
XPCT = 108'b000000111101101110000001011001110011011001111001011010000000101110110110100010001111100001100001000110001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19000

pattern = 95; // 19000
ALLPIS = 207'b110111110110011111001001000100010111010100111010100101010110001001101100001011010100110010110110000110000001001101010010000101110001011100001111100000011111001000110101100000100111010001100110011100100011110;
XPCT = 108'b110100001011101000110011001100100011010111111111011011000000111100101010110001101100101010011111100000100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19200

pattern = 96; // 19200
ALLPIS = 207'b100011000001011010111000011010111110001100110010110100001100110010100100110010101001001111010111101001010101101011111001100000011011001101000111010110000011100101101111010101111111001100011100000100101111011;
XPCT = 108'b111010101111100110001110000000101111011111111100001011111111011011011111001110011111111101100110001111000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19400

pattern = 97; // 19400
ALLPIS = 207'b100101100011001010111001000011010101000110101100001100000110100111000101101111001101100100000011111100101000001000100100110110010000011010010101010110111001001011101110011110001010010010110000101000101011000;
XPCT = 108'b111011110101001001011000010100101011100011111100101111011111011100001111000110001101111010011000010100001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19600

pattern = 98; // 19600
ALLPIS = 207'b101100001101011000010110101010010001011010101010011011011010000011011101000111111010110001111011110110100001111100111111011010001111010111001110000101011000110010010101000010110011110001011101110111110010000;
XPCT = 108'b110000011001111000101110111011110010111101110111111111001111101001001111000110101101111100011001011110111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19800

pattern = 99; // 19800
ALLPIS = 207'b010100011101001000100000101111011001101010010100101000011010001000101000101001110000101101100011111001110010100011011001010110000000011000110001110110010100000111010100010110010111100000010101101100001111010;
XPCT = 108'b000010110011110000001010110100001111101111111001111110011111100010011111111111011011111101000001100101101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20000

pattern = 100; // 20000
ALLPIS = 207'b101011110000011011011100101100111110001010110001111111001100010101110101001001010101000110101000110101110110110010111101011011100110101111100011101011010111110010100000001100011001101010000110010110111111100;
XPCT = 108'b110001100100110101000011001010111111001111101111010001001001101001011110100110110100111111100001101111010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20200

pattern = 101; // 20200
ALLPIS = 207'b000101100010011000010010001110110010011110010010010001011111101101000010101010011011010000010111001001000111010000111001110110011010000110111010101101110111110111011001000101111101000110100011010100011100001;
XPCT = 108'b000000101110100011010001101000011100111101111010101110011001010101001110011100001000110001000000101011101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20400

pattern = 102; // 20400
ALLPIS = 207'b001000101100010011000010010001110110010011110010010010001011111101101000010101010011011010000010111001001000111010000111001110110011010000110111010101101110111110111011001000101111101000110100011010100011100;
XPCT = 108'b001001001111110100011010001110100011110001011000101110001111001011011111101111000111111001000000001111000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20600

pattern = 103; // 20600
ALLPIS = 207'b011010101010110100101011000011000000110000000101010100011100101110001011111010110101101110111011010100010001100101101110100110011110110010011111000100110011001000111111101001100001001100011111101110110110010;
XPCT = 108'b001101001000100110001111110110110110010110111001011010001111011101101111100101100110110011100001000011001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20800

pattern = 104; // 20800
ALLPIS = 207'b110011101001100111011111101010011011100001111110110111010111000111111010001101000110110100100111100010111101001010011010010010001000000011001011001100011101110011111101111001000110011110001010010100111100101;
XPCT = 108'b110111000011001111000101001000111100010111111111011011001111111111011111101100001100110110111001111100000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21000

pattern = 105; // 21000
ALLPIS = 207'b000111001110111110100011010100010110011011101100101100110101111100001111011101110011110101100000010110101111001111110101000011000111101100111100111100000110111100000101000001100011100101110101101001111001111;
XPCT = 108'b000000001001110010111010110101111001010001111001011010001111000101010101011101110010111101100001110100111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21200

pattern = 106; // 21200
ALLPIS = 207'b111011110011110100101000101111101111100111110001110101100101000011111111000001110000001111101000100011010111100010110100000100011101101000010010111000010001011110001000110111011011100000010110001110011110011;
XPCT = 108'b110110110101110000001011000110011110001111111111011011110110001101001011111000101010100101111111110001110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21400

pattern = 107; // 21400
ALLPIS = 207'b000101011110010011001101101010010000001000101100110111100100000110001111011110001111000000010001101111001001111011111010110001010010001101111101011101111000001001010110111000011110011010100000000101111100010;
XPCT = 108'b001111000111001101010000000001111100101110111011111110010000011100001110001010001000100010011111111000110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21600

pattern = 108; // 21600
ALLPIS = 207'b000101001111000110000001010010110011011000001011111000110110100110110001010001110100010110111001110111001010111100101110011111111110100100100111001100011101011001011000100110010110111010000110011001100001011;
XPCT = 108'b000100110011011101000011001101100001101001110000100100011111000011001111100111010001111111100000101010010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21800

pattern = 109; // 21800
ALLPIS = 207'b010101001001000000111001000000110110000111101000110110011011011001001111101100001110111000100110011010001011000000011001110000100100101111100111111010101111010110100001111100110000011001011100100001011101100;
XPCT = 108'b000111101000001100101110010001011101111011111001111110001111100010001111010111100000111010011110000010000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22000

pattern = 110; // 22000
ALLPIS = 207'b101011000010101101110011100011100100110100001100100101001111011010111010111000001111111110111100111101101000010101111110110101100100000111110000110000100100101101000011001111111011010110110001011101111110011;
XPCT = 108'b111001111101101011011000101101111110011101111111010001110000100110001110100000010100100110000110001101111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22200

pattern = 111; // 22200
ALLPIS = 207'b001010110000101011011100111000111001001101000011001001010011110110101110101110000011111111101111001111011010000101011111101101011001000001111100001100001001001011010000110011111110110101101100010111011111100;
XPCT = 108'b000110011111011010110110001011011111001111110011011010001111100111011011110101011000110100100001101000011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22400

pattern = 112; // 22400
ALLPIS = 207'b001011010100011111000011010100111001111000001000101000000001001100011000111000100111010100101011001101011001011001000111001001001100101100100010001010011110111100001010011000111110010011101000010110100001001;
XPCT = 108'b001011001111001001110100001010100001001101111000001010010000011000111110010000000110100000111110100000010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22600

pattern = 113; // 22600
ALLPIS = 207'b100101101010001111100001101010011100111100000100010100000000100110001100011100010011101010010101100110101100101100100011100100100110010110010001000101001111011110000101001100011111001001110100001011010000100;
XPCT = 108'b110001100111100100111010000111010000111001111101111111101001001111010110001101000000111100000001010001101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22800

pattern = 114; // 22800
ALLPIS = 207'b111001011010100011111000011010100111001111000001000101000000001001100011000111000100111010100101011001101011001011001000111001001001100101100100010001010011110111100001010011000111110010011101000010110100001;
XPCT = 108'b110010010011111001001110100010110100110011111111111111111001100011001110101101010000111000000000100111011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23000

pattern = 115; // 23000
ALLPIS = 207'b010011000100000001111100010011101011111110001001000111011111101110111011101100011100010101101011010111100111001001111111011010100111110001101100111011001000010011000000001100101000100010010001110111001100111;
XPCT = 108'b000001101100010001001000111011001100000111111011011010000000000100111010111010111100100000111000111000011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23200

pattern = 116; // 23200
ALLPIS = 207'b111101110011010010000000100111100011100011100101100000110000001010111101011001000110101110111101001000010100011110110001110000101010011101010010011010010110000001101000000111110001010000111001101101111011100;
XPCT = 108'b110000111000101000011100110101111011101111111101111111101111101000011111110111011111111101111001011101101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23400

pattern = 117; // 23400
ALLPIS = 207'b010000100011110111000101001010100011100011000110000100100000000000000101011011001001111011110101110010101010110001001110011011011101010100010001001001100100011000011000110100000000110001100000100000011111101;
XPCT = 108'b000110100000011000110000010000011111100011111001111110001111001101001111110110101010111100011111000010100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23600

pattern = 118; // 23600
ALLPIS = 207'b110001000000011111000100111010111111100010010001110111111011101110111011000111000101011010110101111001110010011111110110101001111100011011001110110010000100110000000011001010001000100100011101110011001111000;
XPCT = 108'b111001010100010010001110111011001111110011010111111111111001000101001110111100110001110011000001111101101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23800

pattern = 119; // 23800
ALLPIS = 207'b011000100000001111100010011101011111110001001000111011111101110111011101100011100010101101011010111100111001001111111011010100111110001101100111011001000010011000000001100101000100010010001110111001100111100;
XPCT = 108'b000100100010001001000111011101100111110011111011111110001111000010100101001111011100111101000000101111011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24000

pattern = 120; // 24000
ALLPIS = 207'b011001100111001111000001110000000000010001011110100111001001100000110101000001111100101101110101001001101100011000010110001101110111010110000110111110011101000101000000011000010011100000101100011001110001010;
XPCT = 108'b000011000001110000010110001101110001101011111011111110011111011110111111100111111010110101111001111001000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24200

pattern = 121; // 24200
ALLPIS = 207'b011101001010110001100001101010001110101011100101000101011010101111100011011010000110100011011001111011011110000000011010010011000101011100001001011011010110101010111101111110111110101110011101010011011001011;
XPCT = 108'b000111111111010111001110101011011001111011111011111110010000101111111100100011100000100010000000000110001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24400

pattern = 122; // 24400
ALLPIS = 207'b101111101110111010101100101000001001101110001100111010100010111110100100100010111110101101110111011011111011101001100000001111100111111001010011010011011001001110110111011000010011010111111101010010100011100;
XPCT = 108'b111011000001101011111110101010100011011011111101011011100000111110011100100010010011100101111111101000001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24600

pattern = 123; // 24600
ALLPIS = 207'b100111000100110001000000111101001100111111111000100110100111100100011101111101101001101101100011101110000011010010011000100101101000101110011101111110101010010011111000101101100100000011011110010100101011100;
XPCT = 108'b110101101010000001101111001000101011000101111100001011101111010111111111010101110000110110100001001101000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24800

pattern = 124; // 24800
ALLPIS = 207'b111000011111011111000010011100111010101001111111011101100001100100111000110111011001011001001110101110111110001001111101101100011101110111011011011110000001110010100011011111110011000000011101100011100010010;
XPCT = 108'b111011111001100000001110110011100010111011111111111111111111010001010101001100000001111111000000100001110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25000

pattern = 125; // 25000
ALLPIS = 207'b100111100110001010110110011101000000001000110000110111101011111000001101100001000101110101000100000110111101100101111001001110100001000101010000100100101001000011100000101000011000011000011010010001111011110;
XPCT = 108'b110101000100001100001101001001111011001001111111011011000000110110101110010000111001101110111110101010000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25200

pattern = 126; // 25200
ALLPIS = 207'b101100001011111110010101101010110011100101001110111101000110000001101001100000000011111010011110010111111100111110011100100101110000110000000111000001110100100010001110111011111101001110100011010110011000001;
XPCT = 108'b111111011110100111010001101010011000101101111110101111101111000011100101010110110000110011011000001010001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25400

pattern = 127; // 25400
ALLPIS = 207'b011001101001110100001010111100010001111010001010100001101100011111110011110111000110101111110011001111101000110010011111001101100000010011101100100101000011010000101100101110010011111010010110101110000101101;
XPCT = 108'b000101110001111101001011010110000101101111111011111110001111011001111111000110010011110100011110100100001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25600

pattern = 128; // 25600
ALLPIS = 207'b111110001101100001101001111010100011010100111111010010010111000100101111111101110110011111000000011100000011110000011110111000111001100100110101001010111001110000010110111100011110100011100011000111010001000;
XPCT = 108'b111111100111010001110001100011010001001110111101011011111111011100011111111111110010111110111000110100110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25800

pattern = 129; // 25800
ALLPIS = 207'b001100110111011000110010101001110100010001011110111010010110011010011100100011111101100000100101100000110010010111110000000111011110100110110100010011000010010010000100101001000011111011101110001000101110100;
XPCT = 108'b000101000001111101110111000100101110100001111001111110011111000000011111111110010110111000111001011010011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26000

pattern = 130; // 26000
ALLPIS = 207'b011110001100010000110010000001011101000010110010100111000111001110011101010001111001000100101110011111100000110111000001001000001110110011010100001010001000001101011111100011011011100000110001101000100111001;
XPCT = 108'b001100010101110000011000110100100111011011111011011010010000010110001110000010011100101110011110000110001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26200

pattern = 131; // 26200
ALLPIS = 207'b111100111001011111000010110001001101011001001011110011011111011100011011111011010110000010010001111000111001101111110111111000111110101101111101001011100100011110011000010011110110110010011100010000000001011;
XPCT = 108'b110010011011011001001110001000000001101011111111111111011111000011001011011100001001111101000001110010000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26400

pattern = 132; // 26400
ALLPIS = 207'b101001001111001101000110000010100010001011010110101000100111101111101001101001001001111111000001011111001111001101011011000001101100111101101110011111000011000110111101111110001011111100110100101001110110100;
XPCT = 108'b110111110101111110011010010101110110110001111100101111101111101101110111110111001000110100111000001001110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26600

pattern = 133; // 26600
ALLPIS = 207'b011110101010101110101101100111011000111000100000101000010000010111000100011100101000001101100011111111001011001011100000101110110000101010111001011101010111110011110110000001101000011000101000100100110100000;
XPCT = 108'b001000001100001100010100010000110100000110111001011010000000000000111110011000001111101010011111101101010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26800

pattern = 134; // 26800
ALLPIS = 207'b001100111001010011101101101001110011111110100100101000001101010010111111010101011110101010111000010101111011011100101101101100110001100011110111101000010110111111110110000110000001100111001100101011011110101;
XPCT = 108'b001000110000110011100110010111011110100010111001110100011111101011011111010111111111110110011000110000011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27000

pattern = 135; // 27000
ALLPIS = 207'b010011100000111011100000101011001100010111111011000110101101010110100001100101000011111101010110011110011001001011010111100101001110110001001001000100010001111001000101101001110010111101101010000101111100011;
XPCT = 108'b000101001001011110110101000001111100011111111001011010010110001101101111111011101010100100011110110000000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27200

pattern = 136; // 27200
ALLPIS = 207'b011001010000001101000100100111101001110110000110110011011110110010011101000101110000010000011010010110100010010000001001111010001101110001111110101110101101110000100000100101011111100100111101010101100111000;
XPCT = 108'b000100100111110010011110101001100111101111011011111110011111000011001111000100000100111101100000111110000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27400

pattern = 137; // 27400
ALLPIS = 207'b101010011001101000001100011001100111001100110010001101100110101101010010010000111100011111111000011110011100111011000011011000011000100111011110011011110101010111001010001101000011001110111000111101011000010;
XPCT = 108'b111001100001100111011100011101011000000111111110001011101111110000001111011111000101110010111000010011101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27600

pattern = 138; // 27600
ALLPIS = 207'b100001100110100100110011111001101110001010010011100011000000101000110111101011111110000111000100001101010000000100100110001100100010110100101111101010101111111011111110001101110001000110011000010001101010100;
XPCT = 108'b111001101000100011001100001001101010101001111110100101000000010101111110010001101000100111111110100100101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27800

pattern = 139; // 27800
ALLPIS = 207'b100101001100010100101100001001100101110101001000001010111011011110011111011001010111011010001101011000100110101111001010011111111011101100100011000101010100111101110101101101011110011010001101101010100111111;
XPCT = 108'b110101100111001101000110110110100111111011110101111111100000000111011100110011111000101110111001111110110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28000

pattern = 140; // 28000
ALLPIS = 207'b000011001110101001111000111001011100000001011011111111001000101001110010111101001101100011001100100111100110011100000111111010110111001100011000010110111111001001101101010110011001111111001111111000000101111;
XPCT = 108'b000010110100111111100111111100000101011011111010000000000000110111001110100000111010100101000000110011101001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28200

pattern = 141; // 28200
ALLPIS = 207'b101001011011010010010001111011001111101000010001100010110100000110110001000001111101011110110001001101111100001001100001101101011001101001011111011110010000010010001000110111010111000100001010001111111101000;
XPCT = 108'b110110110011100010000101000111111101101101111100100101111111110111111111100111100000111110111111110000101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28400

pattern = 142; // 28400
ALLPIS = 207'b010101101010111000010000111001011001001111000000011101010011011010011011111000001001010001011011101011010011010001100000011100010000011001001010001011001011100000110101110101101100100001100110001101010111101;
XPCT = 108'b000110101110010000110011000101010111110111111011111110000110011111001111000001101100101111011110001101011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28600

pattern = 143; // 28600
ALLPIS = 207'b111001101111110010011011000011010110101110110011011101101100110001111001011011001100011101110010110101011000000001101111011111110010100101100110001100110001111000101001110100100100111000100111010110010101000;
XPCT = 108'b110110101010011100010011101010010101110111111111111111111111111010111011000110101111110101011000010111010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28800

pattern = 144; // 28800
ALLPIS = 207'b111011101011100110000000001001111011000111010110101011010000101110011110100101100000100110001010001001011100100011110101100110010101001000010101010011111101011110101011001001101000111111101100111100011110111;
XPCT = 108'b111001001100011111110110011100011110010111111111011011001111000110011101101111100110110110011001010110110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29000

pattern = 145; // 29000
ALLPIS = 207'b111001001001111101001001000100100001001000101001011001010111001100001011000010000011100110111010110011011101100001100111010111011001100100111000010010000110010011001101110001111110101000000101101100000011000;
XPCT = 108'b110110001111010100000010110100000011111111111111111111011111101000101101000110111100110010011000010010110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29200

pattern = 146; // 29200
ALLPIS = 207'b001011010100001110010000000011001011010011010111101011000100101101010010001001010101000110101011110110101100110111001000101000100101101111000000001100011111111001011000000100011100100001010011110010010011000;
XPCT = 108'b000000100110010000101001111010010011001001111010001010011111011000001111110100011010110100000000011010000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29400

pattern = 147; // 29400
ALLPIS = 207'b111000011000101000100001100100111100111100101000000100100000110000010001001100101111000011110001110010100111100001110100001111100000001010111001110100010001011010011110101010011110100010101001100000110100100;
XPCT = 108'b111101010111010001010100110000110100101011111101111111011111111000011111010100100110111110100001100110110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29600

pattern = 148; // 29600
ALLPIS = 207'b000110100101110000011110001111010100011000000010110001110100101011110111100100001010010101011101110111111101101001101111101011010010011110110001110101011111011011111110111110011101110011100000001100000011000;
XPCT = 108'b001111110110111001110000000100000011001111111010000000011111001000110101110111110000111011111110101111010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29800

pattern = 149; // 29800
ALLPIS = 207'b000110100110101100001101111110111110001101110011010111011000000101000011110011010100110101010111111000100000100111101100011011010110110010011011111111011010010110000111011010000100111100111010010001011110011;
XPCT = 108'b001011010010011110011101001001011110010011110011011010000000010101001110101010000001100000011000000000011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30000

pattern = 150; // 30000
ALLPIS = 207'b111010101011100111101011010010010011011100110111001100110000100101110101101100000100001011000110101111010000110100011111101011110011110110000111011011111111010001011000100010100010011000111011001110010111011;
XPCT = 108'b110100011001001100011101100110010111000111011101011011101111111010011111011101111110111001100110111011000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30200

pattern = 151; // 30200
ALLPIS = 207'b010011011110001011100010100011000110100101110100011110100110000000000101001010001100100110001101011000011000110101011010101111000110000111001100011011000001010001001111000000000000100000011000110111011100101;
XPCT = 108'b001000000000010000001100011011011100010111111001011010001111101110000111011111001011110111100001111110101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30400

pattern = 152; // 30400
ALLPIS = 207'b111010110101000100001010011110110110101100111001001001010001111011100100000010001011101011010101001111000001110100001011010111010001000101001011001011110110110011111111001110110000101011110111110110100010000;
XPCT = 108'b111001111000010101111011111010100010011111111111011011101111101000111111101110000101111010111111111000111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30600

pattern = 153; // 30600
ALLPIS = 207'b111110000101011011101100101111011010101011010111111010000100100101010100111000101010100000110001101000000101010110001100100101101010110000001010101011011001011000010111000001100000110011111011011000011100100;
XPCT = 108'b111000001000011001111101101100011100010010111101011011011111000010101111100100011111111101111000010011100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30800

pattern = 154; // 30800
ALLPIS = 207'b101100101100011110110000010100011111101010011000110011110010010111001110111011101011010110100010011000001110111010100000001111001111100101000001101000010110011010110010110101110000011011111011110010010000010;
XPCT = 108'b111110101000001101111101111010010000101001101111111111000000010110001110010001011000101010011000001011010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31000

pattern = 155; // 31000
ALLPIS = 207'b100111010000010111110001101100010101111011110100111110001000101011000001111100010101001110001101001010101000101110100001101001010110010111011110101000001100000111110111000101111101011110000111101111101001100;
XPCT = 108'b111000101110101111000011110111101001011101011101011011101111111110001111001110101100110010100000000000101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31200

pattern = 156; // 31200
ALLPIS = 207'b001100111100110010011011001111100011001001000011011011011110000000110101100100011100010001111000011100001001110001011111010100000011101011000111000100100001001010011010111100110000001101110000011110010001101;
XPCT = 108'b001111101000000110111000001110010001101111111010100100000000110010001010010000110000100100011111001000100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31400

pattern = 157; // 31400
ALLPIS = 207'b100011111100011000111101110001011000011001101000001101101010011100011100010011100011011001010010110110100010000010101101111011011011011001101000110101000101111100100011001101010110110110010100010000110000100;
XPCT = 108'b111001100011011011001010001000110000011011111111011011100110001011111111111011001011100010011111001001011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31600

pattern = 158; // 31600
ALLPIS = 207'b110010011000001110001001001101011110111000110010111101000110101100111000010001011110001010001011000101001111110111111000010100000000011101110000010000111101011001011100100101100010101110000011000010111110000;
XPCT = 108'b110100101001010111000001100010111110000010101111011011111111001010011111011110001100110010000000010010110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31800

pattern = 159; // 31800
ALLPIS = 207'b101000001101000111111000000110011100001110001001001110000100110111001101001111011001010011100011110001010110111110101110001001000110111101101101100010011101000110110101110110010100111101000101100110111000100;
XPCT = 108'b110110110010011110100010110010111000111111000101111111011111000010011011100111001010110000011110100010001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32000

pattern = 160; // 32000
ALLPIS = 207'b101001011101001100101011010100111010000000000010011011010101010010001010101100111000011100001101001000110110001000101010000001110001011001100110011100000111010111100110110110100011010001111010111101001010011;
XPCT = 108'b111110111001101000111101011101001010100111011111111111110110111111111111100011001111100000011111001010001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32200

pattern = 161; // 32200
ALLPIS = 207'b001011010000011011010000001011001011000111000001001000110100111110011111101010110101001011010101011000100011111001110001101100001011111011001100011100000000010001011011000001001011011111111010101110011110000;
XPCT = 108'b001000000101101111111101010110011110010101111000001010011111100110111111010110001011111100100000010101001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32400

pattern = 162; // 32400
ALLPIS = 207'b001100101110110011000100110100010001100100001011111100010111001000011101101001110110000010100110100010001100001110100011110111001100001110110111010100110011010110110000110100011101000100011100111000010110000;
XPCT = 108'b000110100110100010001110011100010110101001111001111110000000011110111110110010111010100111111111110110000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32600

pattern = 163; // 32600
ALLPIS = 207'b011010001110101001111111001111010111011011110001011001111100011011110100110000111101010110010111100010011111000010000110010000100000111001001110100100110010000100011100101100101100011001011010101111111101011;
XPCT = 108'b000101101110001100101101010111111101000110111011011010010000101011011110010001100100101001111111111111111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32800

pattern = 164; // 32800
ALLPIS = 207'b100111010110111001110100001000111111111111011000100110100010101101000101101101000100011100100000001110010110111001100010010001111000110010000100100001001100101001100101010101110100011001110011011101001000011;
XPCT = 108'b110010101010001100111001101101001000011101001101011011110000010101111110011000100011101110011111110000010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33000

pattern = 165; // 33000
ALLPIS = 207'b101000111100010100111110110000100111000100110100111010000001111100100100100111110100000001011010110110100100111010000001011000101000111010010010101100011110101110101111011101010001110001001000011101000010111;
XPCT = 108'b111011100000111000100100001101000010111111111100101111010110101011001111001000010011101100111110100001001001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33200

pattern = 166; // 33200
ALLPIS = 207'b111010110100010010100010111101000011110100100000100000000000011001001111001100010010000011110100100111100100010110110001111001110110101100100011100111101110001000100111001001011100000001001110111100000100011;
XPCT = 108'b111001000110000000100111011100000100011111111101011011001111100100111111101110110111111111100000011100010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33400

pattern = 167; // 33400
ALLPIS = 207'b100001011000000010010101010111001000111101010001110111011110101001010011110001110010011111110100000000011100010100000001001111110111111011110110101111101000110111100101011001111111110011011000111001101001000;
XPCT = 108'b110011001111111001101100011101101001111001111111111111111001000001111110100100100001110011100001000000110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33600

pattern = 168; // 33600
ALLPIS = 207'b011000100000010011100111100101111011101101101011101110101001101111101100100110101000110000111100000110001011000100110001011101010011100101010111001110011100111101011100110111011010010101010010100100111000010;
XPCT = 108'b000110110101001010101001010000111000101111111001111110000110100110101111011010001010100101100111000011001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33800

pattern = 169; // 33800
ALLPIS = 207'b001011001000001111110001101100001001000000110101110011010010010010011000001000010110011000111010100101100101000111001100100011000111011011000111101011101001000001100101110101101111001110010100111101011101111;
XPCT = 108'b000110101111100111001010011101011101010101111011011010000000011101111000101001110100100100011110000001100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34000

pattern = 170; // 34000
ALLPIS = 207'b100010101000000001011010000111001010111010011000101101000000010101001111101111011101101101000100111001111110101011010110010100001011100011001110101111100111000000001011111111111101110001010111000100001111001;
XPCT = 108'b111111111110111000101011100000001111011111111110001011101111101010011111100100110000111100000000001100101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34200

pattern = 171; // 34200
ALLPIS = 207'b101010010010110101011100011001000010000100010000111011000000001101010100100110001110011110001001000101111010110000010010100000110000010100110011001110000000101010110100001011110110011110110110011000001001001;
XPCT = 108'b110001011011001111011011001100001001001011111111011011101111111110111111011100110101110001100000110010000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34400

pattern = 172; // 34400
ALLPIS = 207'b100010010000111010111111000100011100111011001000100110000001101110010001000110101000010110111110010100010100111100110000001011111111001111111011100100001011100000000011010101101001010001110111100100000111101;
XPCT = 108'b111010101100101000111011110000000111010111111101011011001111111101101111100100001011111101100001011001010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34600

pattern = 173; // 34600
ALLPIS = 207'b011011110100000001110100111110001001100111111000010101101001010111110011010101010101001011110011100011011010110101001110101101110001100011101110001011101101100001101001010100100100011001111000010001110010001;
XPCT = 108'b000010101010001100111100001001110010010011111011011010011111100111011111011100110111111111000001101001111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34800

pattern = 174; // 34800
ALLPIS = 207'b100111011110010001001111101111000101101001001110010111010101010111011111011100110001100110110010101000111100110100111011111100101001110001111110010001111001010101011101010111000011010100011110001000001001100;
XPCT = 108'b110010110001101010001111000100001001010011111110001011001001011100111110110101010000111000100000001000010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35000

pattern = 175; // 35000
ALLPIS = 207'b100111001000001010111101001001110010010100000101011101010011111111011110111000100011110011111100100110001110011011011100011101010011000011000000100111011000011001011101111001111001010011000110011100101110111;
XPCT = 108'b110111001100101001100011001100101110011111111110001011000110000110001111101010011100101111011110010101101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35200

pattern = 176; // 35200
ALLPIS = 207'b110011000011011000110111100011110000010100110001001101011111000000101001100000100110000111110011001111110101100110000000011100000110010110000011110010101000011111101111111000011100001011100000010000000001011;
XPCT = 108'b111111000110000101110000001000000001011011111111011011011111110110011111101100101000111110111000001011101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35400

pattern = 177; // 35400
ALLPIS = 207'b000001001110011101001110011101001010010000110001110111110011000001001111111000010110101011110000111010011000010110010101011010110100110111011110001110101111110110100011011000001101011100000110110011111101000;
XPCT = 108'b001011000110101110000011011011111101110011111011111110010000110100011110010010111110100010111111111110011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35600

pattern = 178; // 35600
ALLPIS = 207'b010010111111000010110000110100110000100100010000111111101111101001100010110111111001001110111011001110000101100001000101010001011011001100110011011010001110001011101010000110110010101100110001010001100100000;
XPCT = 108'b001000111001010110011000101001100100001011111011011010011111101111111111011101001101110010111110000000111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35800

pattern = 179; // 35800
ALLPIS = 207'b101110000000000001010111110110111110001101001110101100010111011100000001111101100000000001010001111110001000111110001001111010010101000100110100111010101011100000110011100101110010010101100001010111100101000;
XPCT = 108'b111100101001001010110000101011100101011101111101011011000000111000011110101011011110100101011111110010110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36000

pattern = 180; // 36000
ALLPIS = 207'b000011111110001001000010110011100000100001111100011011101010000111000001010010000111101100010100110100101011011101101101111010011100000010111001101011001010111100001101000101111001011100000100010110000111111;
XPCT = 108'b000000101100101110000010001010000111011101111010001010000000010000111100000011011000101001011111010100000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36200

pattern = 181; // 36200
ALLPIS = 207'b111101100101001111010011111000010110011010011101000110100000001001100110010010111110101100100011100110111011011000010001011010100010000101111000000110101000000110001001000000000000000011101101111111000100110;
XPCT = 108'b110000000000000001110110111111000100110111111101111111101001100100011110110101011111110000111000010111001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36400

pattern = 182; // 36400
ALLPIS = 207'b001101111000110110010101000001001011001001100010100000010001100000011000011101100100000000010101110000011101100000110000111001010000111001001110101001010000100011000100000000111000000011011110111000011010001;
XPCT = 108'b000000001100000001101111011100011010101001111001111110011001010001001110000100110000110000000000001010111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36600

pattern = 183; // 36600
ALLPIS = 207'b101111111101000110010110010001011001010101000011111000011100111001010000111001100110100011010110100010011000110011010000100111100001010101100001000100011110010101000100100000110110000001011110001100011001001;
XPCT = 108'b110100001011000000101111000100011001001101111101011011011111011001111111111111111110111111111001011101000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36800

pattern = 184; // 36800
ALLPIS = 207'b110001000111001001011001010000001010110110110001011101111111001100100001000001101101010100100011001011111100000001010101001111110010111001011100011010111001101000110010100100001100011001111100011010101010010;
XPCT = 108'b111100100110001100111110001110101010100011111111111111011111100011011111111110010010110000011000101110000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37000

pattern = 185; // 37000
ALLPIS = 207'b010110010010011110000001011100100101010010111000110011001010010101001101110101010110111100100100110111110110101010001111111101111000011110110101100110100000011101010111100111000110010011000001101010111010110;
XPCT = 108'b001100110011001001100000110110111010010011111011011010010110100111110101000010011100101101000111101111100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37200

pattern = 186; // 37200
ALLPIS = 207'b100101110010010100101011000000111101000000001011100100000110111010111011100001110001010100001101110001111001110101101011101010111011110010100000111110111011101100000111100010001000001100011001111101011111101;
XPCT = 108'b111100010100000110001100111101011111110111110101110101001111011000001111110111111000111010100000011010001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37400

pattern = 187; // 37400
ALLPIS = 207'b101110110000000010011111001000101010111100001100110100000000000110100110000101110011001110100000101111100000011000001101010011110110010100110101000001111000100001001001101000101000000000001100100111000110000;
XPCT = 108'b110101001100000000000110010011000110010111111100001011110000100110011110100011110110101111111111110100101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37600

pattern = 188; // 37600
ALLPIS = 207'b011110111100100110000010010010111001010000001010010110010001101110100010000110100000100111110110101011110010001000100001111100110010001110000101110100100001001001101100111110011110010000111001111001100110011;
XPCT = 108'b000111110111001000011100111101100110001011111001011010000000100000001010110010000010101101000000000000001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37800

pattern = 189; // 37800
ALLPIS = 207'b100001111000110010111110010010111001101010101000010101101000101101010000000000100001100000111010011010110111100100110000110001010001100101101111010100100000011101010101110000100011000001110011000001100111001;
XPCT = 108'b110110001001100000111001100001100111110011111111111111010110100111101111100001001111100001011111110111001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38000

pattern = 190; // 38000
ALLPIS = 207'b011101001100111100010001110111110000010100101010010100101010111110001011011000011100101010110111001000100001010011100111100010001111000000111000111101010101100010100100000101010100000000010010010110001001010;
XPCT = 108'b000000100010000000001001001010001001101111111001111110010110111111001111101000010000100000111111011101011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38200

pattern = 191; // 38200
ALLPIS = 207'b001111100110000111100101001010001011001100011000111000001011110010101101101100111111101101001000101101101100101101011110101111010111101100110001011100001111110011010010000100000100100000011000000000010111000;
XPCT = 108'b001000100010010000001100000000010111000001111001011010010000110011101100010001011111101111011110100011110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38400

pattern = 192; // 38400
ALLPIS = 207'b101011010110010011101011011110001000011001101111011000111011000110010101110011010110001111111110001010110000101111110101111110001011011000110000100000110001111111111110111110011100001010111111011110101111001;
XPCT = 108'b111111110110000101011111101110101111001111111100001011110110111110111111001000100110101001011111010001001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38600

pattern = 193; // 38600
ALLPIS = 207'b110010100100011010001010100000011101100001010000010110000001101100001111001101100000011000110001011011111111011111010100111011101110011011110011011111000100101001101111010100000100010111110111010110010000000;
XPCT = 108'b111010100010001011111011101010010000010111110101011011101111000000010101000111011011110101100000100001000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38800

pattern = 194; // 38800
ALLPIS = 207'b111100011110110110110000000011011101100100010010111010100010001110000011001100101101101010011001101101111111111011111011001010010100010001100010001111000000000110101110000000111101001101110101001100101110010;
XPCT = 108'b111000001110100110111010100100101110101111101101111111110000111100111110111001101111100011111110010100000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39000

pattern = 195; // 39000
ALLPIS = 207'b101101111010000011011000101001111000100101010111110011000100100011000101010011111100110110011111001011001011011101101001011000010001101000101001110101000111111000111101000011011111101001111100100110010110000;
XPCT = 108'b110000010111110100111110010010010110111111110110101111010000100010101100100001001101101010011111100000010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39200

pattern = 196; // 39200
ALLPIS = 207'b110101100100111101110100011011010110101110001100001101110100111101001010010110010010111101010101000101010111111110000111010001111010000110110000110001000011100001010100010101110110110010101101101111100001010;
XPCT = 108'b110010101011011001010110110111100001101111101111111111110110001101111111000010110101100101111111001101001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39400

pattern = 197; // 39400
ALLPIS = 207'b011010101101110110111000000111100100101101001010111000011111101001000111001110111110010101010101111100011101001010111111101001001001011011111001101111101001100100101101000111010111011100100110000001101110011;
XPCT = 108'b000000110011101110010011000001101110011011111001011010001111110011111011100111001111110000100000000011101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39600

pattern = 198; // 39600
ALLPIS = 207'b100011111010011100100000011010011110010110011100110110100111101100001010100000001111101100001110010100010100101101100101101101111010110000010100100001101110000101010011000111001100100100011101010110100110100;
XPCT = 108'b111000110110010010001110101010100110010101111101011011101111011111011111111110110000110111000001011101100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39800

pattern = 199; // 39800
ALLPIS = 207'b111101100110101111110001100111101010001110010101101111111000011111100101101010101010000011110011001110111110111101100100000101010100001010101010101110001110000111011101010111111110111011100000111100100110110;
XPCT = 108'b110010111111011101110000011100100110111111101111111111000000011011001110000010111001101000100001001010011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40000

pattern = 200; // 40000
ALLPIS = 207'b011100000000110001001111101110111000010010011111110111111111100101011100001010010100110101000011111101000000010101010010010010010101001001010101111010000010110110000001111001110111110010101010110011011001100;
XPCT = 108'b000111001011111001010101011011011001111011111011111110010110001100001111000001100000101100011110111011011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40200

pattern = 201; // 40200
ALLPIS = 207'b000111111000001111110110110110000010000000011011011110011001110100010101111110100100011010000110000001100011101000011100111100100111001000000101111110010101010100100111000000011100001001100010011100111000110;
XPCT = 108'b001000000110000100110001001100111000011101111001011010000000001111001110011000011111100110011110001011000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40400

pattern = 202; // 40400
ALLPIS = 207'b010001011010011100111110011100010010111000110010110111011010101011000010101110000111110110100001101110011011010001010000001011111010010001110111110001110000001100111100100001100110101110000011101000001010101;
XPCT = 108'b000100001011010111000001110100001010100011111011111110001111110010011111111100010011111011100000000101000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40600

pattern = 203; // 40600
ALLPIS = 207'b000100001010110000011011110000000000000101100000001011110101111111111111100001101011111100001101111100101001101111111110010100011001011111111101010000001111010010001100000101101111010101001001011110010100000;
XPCT = 108'b000000101111101010100100101110010100100111111010100100011111010011011111010100001101110101100001011111011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40800

pattern = 204; // 40800
ALLPIS = 207'b111111011000100100111010000110100101001101001101111110010110000011101110000100101000010000101000110110001011101011001111110110001101010111001010100000101000111010101001010101011111010110100010111111110011001;
XPCT = 108'b110010100111101011010001011111110011011111111101011011010000100001101110000000001011100101111110000110110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41000

pattern = 205; // 41000
ALLPIS = 207'b011000010010011011000011100011100100100010010100101110110011100100000100110010101100010010001010111010111000110100100011110100011100111001001011011111110111010110010111011101101010111100110010101011110111111;
XPCT = 108'b001011101101011110011001010111110111110011111001111110000110011101110101000001000011100000011111010101001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41200

pattern = 206; // 41200
ALLPIS = 207'b100101100101010100100111111111011101010001110000010100001101001010000010111111011111000100100100100010010101011110011000010101011001111110101101001110111010100110110010010010111111000111010000000101110010100;
XPCT = 108'b111010011111100011101000000001110010101100111101111111001111010010101011011100000110110101011110000000010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41400

pattern = 207; // 41400
ALLPIS = 207'b100001011000010000001100010110011110111110000101001011111010011010011110111010000000011010110110100101111111111001111001000100001001111110101011000100110101000111001001010111111110100110001110000010000011101;
XPCT = 108'b110010111111010011000111000010000011111011101110101111101001101100101110010110010011111110100000011000000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41600

pattern = 208; // 41600
ALLPIS = 207'b010110011000100111110000110011000101000000110000111011000001000101100110010010101111111111010000101100110110001011111111011001010010011111110111101111011110010010101010000001011001010011000010011001110010100;
XPCT = 108'b001000000100101001100001001101110010001011111011011010001001101111001110111111111101111100100000100011101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41800

pattern = 209; // 41800
ALLPIS = 207'b110111111010001001110010001001001011010011111001111110011001100110100011111110101101000111100110001000111100010010101000111000110001000011111111011100001111110011011001011000001000110001110000111110101001001;
XPCT = 108'b110011000100011000111000011110101001010111111101011011011001111100101110111111000010110111000000111010011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 42000

pattern = 210; // 42000
ALLPIS = 207'b111110100010011100000001011110001011011110011111101101111110110001110000001001010110101111100101101001100010110000001100100101011000100010000001110101111101100011110111011100001101001101001111011100011011101;
XPCT = 108'b111011100110100110100111101100011011010111111111011011110000011111011110101001000001100011111110000100010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 42200

pattern = 211; // 42200
ALLPIS = 207'b110110100110001010010111000001110011011100101000010010000000110000110100011101111010000111000100101010011110011110110110100010001111001111000110110110000101001000101001110000011011011101000010010100000111100;
XPCT = 108'b110110000101101110100001001000000111011111111101011011011001101101111110000110111010110000100001001110101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 42400

pattern = 212; // 42400
ALLPIS = 207'b010100110000110001011010110001110101101110100000010101000000110000001101011110101000010011000111000010010010001011000110110011111000000111100101101111100100000100110110110001101110110101000101011000001111011;
XPCT = 108'b001110001111011010100010101100001111100011111011111110011111110111011111111101111000110100000000010100101001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 42600

pattern = 213; // 42600
ALLPIS = 207'b100010010011111010011001111110110011000001100110011011100010111110000010101101011100101111110110001110011111110101000100100011101001011110100010001001101001110101000000010111111001010110000010010111110010111;
XPCT = 108'b110010111100101011000001001011110010001111101111011011111111101011011111111111101001110100100001111110000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 42800

pattern = 214; // 42800
ALLPIS = 207'b101111000010011010101100110101011100000001010000101100110001100101010110110110010000111100100011011100110110001010011110000100000100100010011100011011001111111000110010011000100001110000000100011101111001101;
XPCT = 108'b111011001000111000000010001101111001000111111101011011100000000001110110110001110011101100011111101011110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 43000

pattern = 215; // 43000
ALLPIS = 207'b011111101100100001000011100011001010011000001010011010001011110111010110011101011111000010110000001010001011001111100111111010110101011101000101100100101010010101101011101110000001101101110110101111100111111;
XPCT = 108'b001101110000110110111011010111100111010111111001011010000000101000111110000011110110100010100001100011101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 43200

pattern = 216; // 43200
ALLPIS = 207'b001111011010011101101110101010000110011010110010100110100010110111010011010000001010110110001111100111101010101011010001010110101010011000011100000111110010101110010000000101010010010010001010111101111001000;
XPCT = 108'b000000100001001001000101011101111001001111111001011010010000100111011010011011011111101101111111000011010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 43400

pattern = 217; // 43400
ALLPIS = 207'b001111111011100010011011011110110001001010101010111101000110011000001010111011100000100001111110110011101101100010011111110100110111111011000100011101011010101000010001011101011100101111110101010011111001011;
XPCT = 108'b000011100110010111111010101011111001011010111011011010011111110011111111100111000001110010100111101011111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 43600

pattern = 218; // 43600
ALLPIS = 207'b010001111010000000100100000000000011001110111101001001001001011111001100110010010010010011010111111110001110101010101100001000011000010100010010110101010101011101001111001001000001111111100000001110000101101;
XPCT = 108'b001001000000111111110000000110000101110111111011111110000110110001011111001010100110101001111110011000111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 43800

pattern = 219; // 43800
ALLPIS = 207'b100001111000000011000001100011100011010010100110010111001110100100110011100110100110100111111010010001010110000010110011000011110110001010100010000110110011101101110101111101010011001010000101000110000000010;
XPCT = 108'b110111100001100101000010100010000000111101111111110101010000010011001110111010011010100101111000100100001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 44000

pattern = 220; // 44000
ALLPIS = 207'b001001111001100010001110110100110000110011110100000101010110100000100001011000000010110110011000001011111100111011100111011110100111000100101101011110110110111001111011100010111111010011010001010001000000011;
XPCT = 108'b001100011111101001101000101001000000111011111010101110011001011000011010001100111110111101100001100010100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 44200

pattern = 221; // 44200
ALLPIS = 207'b010101011000101100111100011110110111110100110010101111100010110111000101101000111101011010011100000001111001000010110110101010100000110100100010100011100101111010010000011000010011111011001010101001101101001;
XPCT = 108'b000011000001111101100101010101101101101011111011111110010000010100101110100000000100101100011111101111000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 44400

pattern = 222; // 44400
ALLPIS = 207'b110101110001101101011010110011100000101100011111111011110100101101111011101110010000010011110111101001010101001110101110101111101010100101101001011000010111111101010011101100011010111011010110110101110101000;
XPCT = 108'b111101100101011101101011011001110101111111110111111111011111001000101111101110101011110001011001010101011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 44600

pattern = 223; // 44600
ALLPIS = 207'b110011100110101100110111100111011111000011101010101011101101111001010111001100100001001011011011111011000010111101011010111111100100111001110000010011101111101000111011101111111001000101110011110101011010001;
XPCT = 108'b111101111100100010111001111001011010011111111111011011110110010011111011110001111011101001011111000101111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 44800

pattern = 224; // 44800
ALLPIS = 207'b001000000111100110110000001001111111010110001011110000010011110010111011111111111001100010110001011010000110101000011010111011100101101001110000101011101111001100110101011010000101100011111100100100011001000;
XPCT = 108'b000011010010110001111110010000011001110101111001110100011111000011011011101101000011111110111111001010101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 45000

pattern = 225; // 45000
ALLPIS = 207'b000100001001110111100111100110010100011110011111101101101000010001100100110111000111011101001101000010110111111100001110101000000110110110111100001101011110010001110110000110110010001111001001010010110101100;
XPCT = 108'b001000111001000111100100101010110101101000000011111110001111110111100101110101001101110011011110100100111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 45200

pattern = 226; // 45200
ALLPIS = 207'b010111001000001100110101101000001000101001000011101010101011000000110011011101001011001100011010011100111011010101110110010100001101101001001001001001100100101010011000010101001011000000001000010001101110111;
XPCT = 108'b000010100101100000000100001001101110000011111001011010000000011010100100011011100000100011011110011110100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 45400

pattern = 227; // 45400
ALLPIS = 207'b110011101110000110011100101011010101001010110100100000101010110011011011000101000000101101011101011101100101111011001001001101000011001001000101010000010111001100011111001100101011111000001001011110010011001;
XPCT = 108'b111001101101111100000100101110010011010111111101011011110110011100101111100000101011101100111110110100010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 45600

pattern = 228; // 45600
ALLPIS = 207'b001101011110011011000001000001101001001000010010001000000100100101101010000000110111110111000011101000101011110001011010010110001101011010010101111111010000110111001010000010001100000011000100111010011111100;
XPCT = 108'b001000010110000001100010011110011111100001111000101110001001111101101110100100110000110000100000101100001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 45800

pattern = 229; // 45800
ALLPIS = 207'b011000000000100010101111110110101111101100011110101100111011001010100110010110000111110110010010001011100001001111101101011011100010010111001010011101111100010100011010100100110100100100010010001010001101100;
XPCT = 108'b001100101010010010001001000110001101101010111001111110011111111010001111011101101110110110000000100010111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 46000

pattern = 230; // 46000
ALLPIS = 207'b111100001111000110110000000011011011100110011100011011101101100010010101000001110101101000011111000100100011101011001110000011011010001101110011001110110001011111111101101001001001000110011011111010110100110;
XPCT = 108'b110101000100100011001101111110110100110011111111111111101111001100111011001110100100110111111000101110001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 46200

pattern = 231; // 46200
ALLPIS = 207'b101001101000010010110111110101110011100000100101001111000100101000110000001101010011100001110000001000000001110010110110010001011101111110010010110100001001100010110111011011100100010000101111101011100100001;
XPCT = 108'b111011011010001000010111110111100100110001111111110101010000010011101110101000011011100011111111100100010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 46400

pattern = 232; // 46400
ALLPIS = 207'b001000101101111110011110000010101011011010100000001011000001001010111001101000010111101011110000111101001110011101001001000000001001110001110101101001011100011011110001001100100000111100001111011100100110010;
XPCT = 108'b000001101000011110000111101100100110110111111011110100001111000101111111100111100101110000011001000000010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 46600

pattern = 233; // 46600
ALLPIS = 207'b111001010010001001010101101000111001000111000001000010011010111111100111110101011010101001011110000001101100010111111001000110100010110111001111000000010110010110011110111100100100111011100010110010011111000;
XPCT = 108'b111111101010011101110001011010011111100011011101111111110000010011001110100001111111101110011110111110001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 46800

pattern = 234; // 46800
ALLPIS = 207'b110100110100001111111110000111110110001001111111001011011110011000011100101000010000101000010100000001110101000011001001111011100000100111001110001000101010010110101111111001010101100110001010111001100111101;
XPCT = 108'b111111000010110011000101011101100111111011111111111111101111101000111111001100110000110110000000111000011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 47000

pattern = 235; // 47000
ALLPIS = 207'b111111100100110111100011001011100000100111110101010110110100011001111000000111000010101010111011100010101101100010011011010101011101001000101011010001010110011000001100000010110100000010100110010010111111100;
XPCT = 108'b110000011010000001010011001010111111001011111101011011100000111111111000010011111111101111011110100110110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 47200

pattern = 236; // 47200
ALLPIS = 207'b101010110100110101111111100011000100100101011000110010000001111100000110010101000000100100101011100100111100111100110110110000000100101101001101010101101110100100010101010001111111000110001000100000101011100;
XPCT = 108'b110010001111100011000100010000101011011011111101011011011111101000001111101110011011110110100000010000100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 47400

pattern = 237; // 47400
ALLPIS = 207'b101000010000111010101101101001110100011011011000110110100010110010110011101000110001011101110110111000011110111001010000110101111011110001111001101100010111101100100001101111110000111100101000111000001001110;
XPCT = 108'b110101111000011110010100011100001001111011101101110101110000010111101110100010010110100000000111010111100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 47600

pattern = 238; // 47600
ALLPIS = 207'b011111100111010011111010010101100111010011011110011010100100010000110000000011010011000110100111001010011010001011101011111111111101000011011100000101101101000110111100101101111010101010011111110111010111001;
XPCT = 108'b000101101101010101001111111011010111001111111001011010011111011101001111010111010110111010111001001000101101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 47800

pattern = 239; // 47800
ALLPIS = 207'b111100001101001010001000110010001110101000000010111100010110001110011010011000111000001101100100111011100000100101000000111111101010110011111011001011011001100001110000011100111011101100001001001001101111011;
XPCT = 108'b110011101101110110000100100101101111101011111101111111111001110010111110010101100011110010000111001001101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 48000

pattern = 240; // 48000
ALLPIS = 207'b101000100000000100101111011110011101101100111101101100000100001011110010101001111000110110000111111111011001110111001111101100001001101011101011000101101101001110110101011001110000010001111111011100110110000;
XPCT = 108'b110011001000001000111111101100110110111111110101110101001111010011111111101101110011111101000001000110101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 48200

pattern = 241; // 48200
ALLPIS = 207'b100110001011100111100101001111011110000100011100011100001000011000010011111011011111000010001010010101111001100011010000110111101010101011011000010111010101101001001111000001000011101110100000000001100101010;
XPCT = 108'b111000000001110111010000000001100101010001111100001011001111000010001111100111101111110001111110001001101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 48400

pattern = 242; // 48400
ALLPIS = 207'b010000001011011110010011001001011111010000110111000001001110011110110000110101000100010110011000111111100010100100101100000100000000111001110000101001000100111010101111000010010011001110101100011101011110101;
XPCT = 108'b001000010001100111010110001101011110111111111011111110001111010011011111001111001101110010111110001011000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 48600

pattern = 243; // 48600
ALLPIS = 207'b011101011010111100110010000111011011100100001000001011101110111110010000001000100001101100000001101111111010011100010111101110100111101111001101100010111011110000111100011100001110000011010010111111101000011;
XPCT = 108'b000011100111000001101001011111101000100111111011111110010000110100011110111010100001101111011001011010000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 48800

pattern = 244; // 48800
ALLPIS = 207'b011101000111100111010100101011001101001010110011101101011001100101101100010011110110101111100111110000101000111101101110010110000011110101101100011100110011001101110011110000001101000000100000110101110110010;
XPCT = 108'b001110000110100000010000011001110110110111111011111110011001101100001110101110101000111111011001110101001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 49000

pattern = 245; // 49000
ALLPIS = 207'b001101001111001000110111101111110010011101001110001101011100000001111110110101100000100001011010000111111111110010110000001001110110011110110111110000111101101010010001000010101110000110001010110011001000101;
XPCT = 108'b000000011111000011000101011011001000110000001011110100001111011010010001001110011101110111111001100110101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 49200

pattern = 246; // 49200
ALLPIS = 207'b111110100010011010110011001110011111101011101111011010111110110001000011000011101101110111111100101001011001111101001111111001001000011010110000101001101011001100101011001111100001011011111110000101001010001;
XPCT = 108'b111001111000101101111111000001001010010111111101011011000000110011111110100010010111101001111111000110000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 49400

pattern = 247; // 49400
ALLPIS = 207'b001001110100101011101001101010010011010111100110000001101111110101001011011011101110000100010110110100100001010010110100101000101101100111101011100101111111001111000011000101010100101101011010101001101101101;
XPCT = 108'b001000100010010110101101010101101101111011111011111110001001100101110110000111001100110001100001111001001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 49600

pattern = 248; // 49600
ALLPIS = 207'b001100111001100101110111110001110000011111010111001110111010011001010001011011100001011001111111010001000111111100111000111001001010101111100111111110110000110011111101000110100011101011101000110101111110011;
XPCT = 108'b000000111001110101110100011001111110110100100000101110010110100111010001001001101111101010111110110010011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 49800

pattern = 249; // 49800
ALLPIS = 207'b001100010010101000110101101101111000100010001111010100111110011001110111101111000100101111000011001110010111110010111110010001111111010100001000010011100001000101011001110011001111010010011000010011000111001;
XPCT = 108'b000110010111101001001100001011000111110001101000100100000110110000001111001001001010101101111111011101111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 50000

pattern = 250; // 50000
ALLPIS = 207'b101110010010010010011000110101100011101010001010101011011001011000100100010110001110010001010011110111000101100111111110001010110100010101111111110110010110111101011001110000110000100001011111110010010111000;
XPCT = 108'b110110001000010000101111111010010111011010010110001011000000101100000000001000001000101111011111100101010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 50200

pattern = 251; // 50200
ALLPIS = 207'b010010100000111011100011100011000100011010100000100010000001010110101011011100001100001001101000010110000101101010010111101000110111001001001111000101010000011000011111100010000000011011011011000110000101100;
XPCT = 108'b001100010000001101101101100010000101010110111001011010001001011000111110100111011110111001000000111111010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 50400

pattern = 252; // 50400
ALLPIS = 207'b101100110111111011111100110100010000100011010010111010001100011011011110010110001111011010000101001100010111110100001001101000011010111111110100110100000101110011101110101011110110010011000110110101000010101;
XPCT = 108'b111101011011001001100011011001000010101111000100101111101111011001100001011111100110111101111001100111111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 50600

pattern = 253; // 50600
ALLPIS = 207'b101010000011101100010111000011101111010011011001000000011000110111111001010011110100101011101001110000010101110000111100100101110110101010001011000010011000010101000010001001111010111011101001100100001101000;
XPCT = 108'b111001001101011101110100110000001101001101111101010001111111101000001111110110000111111000011111000001001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 50800

pattern = 254; // 50800
ALLPIS = 207'b011100001010000010110011101101100111110111010100000101110101001010001000010100011011010100101011111010100111111100001101001100001010011111011101110111111110011101110010000111101011111011010101111000110110101;
XPCT = 108'b001000111101111101101010111100110110100010000011111110010000011010110000011001111101001000111110111001011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 51000

pattern = 255; // 51000
ALLPIS = 207'b101110010010100111011101001111010110100101110000011011101100001100111100011101010100111011011100010011111011010101100001011110000101011100101001001101011000101001001010010101101001111011110110000001101010001;
XPCT = 108'b111010101100111101111011000001101010000011111110000001110000111000101110011011001001101000011110001100000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 51200

pattern = 256; // 51200
ALLPIS = 207'b101010000001011101101001001011001111101000100010111101101110101001111110010001001110011101011001111001110001001110010010100101000111111001101011111110011111000011001100011100011010011010000010011011010011001;
XPCT = 108'b110011100101001101000001001111010011001011111110000001111111111111111111110101110001111001111110011000011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 51400

pattern = 257; // 51400
ALLPIS = 207'b001101101100010011010000100110010110110010100001010110101001000001100101110110101100110110110111000111100111111101101111001111011011010110110111100010010111101100110101001011010011101001100100110101111011101;
XPCT = 108'b000001010001110100110010011001111011111100000001111110000000001100101000100001110111101010111110011000010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 51600

pattern = 258; // 51600
ALLPIS = 207'b110000011110100110101000000011101101110100101000010111000001100100100001011000110101000011001100111011000111111010001100001000100010001001101110011101000110101110101110001000011110111100110010111101001001101;
XPCT = 108'b111001000111011110011001011101001001101111101111111111011001100011111110110100100101110000000001111010110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 51800

      $display("// %t : Simulation of %0d patterns completed with %0d errors\n", $time, pattern+1, nofails);
      if (verbose >=2) $finish(2);
      /* else */ $finish(0);
   end
endmodule
