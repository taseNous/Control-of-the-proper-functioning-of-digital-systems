// Verilog pattern output written by  TetraMAX (TM)  B-2008.09-SP2-i081128_181834 
// Date: Wed Jul  6 12:10:47 2011
// Module tested: c7552

//     Uncollapsed Stuck Fault Summary Report
// -----------------------------------------------
// fault class                     code   #faults
// ------------------------------  ----  ---------
// Detected                         DT       6775
// Possibly detected                PT          0
// Undetectable                     UD          0
// ATPG untestable                  AU          0
// Not detected                     ND        113
// -----------------------------------------------
// total faults                              6888
// test coverage                            98.36%
// -----------------------------------------------
// 
//            Pattern Summary Report
// -----------------------------------------------
// #internal patterns                         208
//     #basic_scan patterns                   208
// -----------------------------------------------
// 
// There are no rule fails
// There are no clocks
// There are no constraint ports
// There are no equivalent pins
// There are no net connections

`timescale 1 ns / 1 ns

//
// --- NOTE: Remove the comment to define 'tmax_iddq' to activate processing of IDDQ events
//     Or use '+define+tmax_iddq' on the verilog compile line
//
//`define tmax_iddq

module AAA_tmax_testbench_1_16 ;
   parameter NAMELENGTH = 200; // max length of names reported in fails
   integer nofails, bit, pattern, lastpattern;
   integer error_banner; // flag for tracking displayed error banner
   integer loads;        // number of load_unloads for current pattern
   integer patm1;        // pattern - 1
   integer patp1;        // pattern + lastpattern
   integer prev_pat;     // previous pattern number
   integer report_interval; // report pattern progress every Nth pattern
   integer verbose;      // message verbosity level
   parameter NINPUTS = 207, NOUTPUTS = 108;
   wire [0:NOUTPUTS-1] PO; reg [0:NOUTPUTS-1] ALLPOS, XPCT, MASK;
   reg [0:NINPUTS-1] PI, ALLPIS;
   reg [0:8*(NAMELENGTH-1)] POnames [0:NOUTPUTS-1];
   event IDDQ;

   wire N1;
   wire N5;
   wire N9;
   wire N12;
   wire N15;
   wire N18;
   wire N23;
   wire N26;
   wire N29;
   wire N32;
   wire N35;
   wire N38;
   wire N41;
   wire N44;
   wire N47;
   wire N50;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N69;
   wire N70;
   wire N73;
   wire N74;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N82;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N94;
   wire N97;
   wire N100;
   wire N103;
   wire N106;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N118;
   wire N121;
   wire N124;
   wire N127;
   wire N130;
   wire N133;
   wire N134;
   wire N135;
   wire N138;
   wire N141;
   wire N144;
   wire N147;
   wire N150;
   wire N151;
   wire N152;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N178;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire N185;
   wire N186;
   wire N187;
   wire N188;
   wire N189;
   wire N190;
   wire N191;
   wire N192;
   wire N193;
   wire N194;
   wire N195;
   wire N196;
   wire N197;
   wire N198;
   wire N199;
   wire N200;
   wire N201;
   wire N202;
   wire N203;
   wire N204;
   wire N205;
   wire N206;
   wire N207;
   wire N208;
   wire N209;
   wire N210;
   wire N211;
   wire N212;
   wire N213;
   wire N214;
   wire N215;
   wire N216;
   wire N217;
   wire N218;
   wire N219;
   wire N220;
   wire N221;
   wire N222;
   wire N223;
   wire N224;
   wire N225;
   wire N226;
   wire N227;
   wire N228;
   wire N229;
   wire N230;
   wire N231;
   wire N232;
   wire N233;
   wire N234;
   wire N235;
   wire N236;
   wire N237;
   wire N238;
   wire N239;
   wire N240;
   wire N242;
   wire N245;
   wire N248;
   wire N251;
   wire N254;
   wire N257;
   wire N260;
   wire N263;
   wire N267;
   wire N271;
   wire N274;
   wire N277;
   wire N280;
   wire N283;
   wire N286;
   wire N289;
   wire N293;
   wire N296;
   wire N299;
   wire N303;
   wire N307;
   wire N310;
   wire N313;
   wire N316;
   wire N319;
   wire N322;
   wire N325;
   wire N328;
   wire N331;
   wire N334;
   wire N337;
   wire N340;
   wire N343;
   wire N346;
   wire N349;
   wire N352;
   wire N355;
   wire N358;
   wire N361;
   wire N364;
   wire N367;
   wire N382;
   wire N241_I;
   wire N387;
   wire N388;
   wire N478;
   wire N482;
   wire N484;
   wire N486;
   wire N489;
   wire N492;
   wire N501;
   wire N505;
   wire N507;
   wire N509;
   wire N511;
   wire N513;
   wire N515;
   wire N517;
   wire N519;
   wire N535;
   wire N537;
   wire N539;
   wire N541;
   wire N543;
   wire N545;
   wire N547;
   wire N549;
   wire N551;
   wire N553;
   wire N556;
   wire N559;
   wire N561;
   wire N563;
   wire N565;
   wire N567;
   wire N569;
   wire N571;
   wire N573;
   wire N582;
   wire N643;
   wire N707;
   wire N813;
   wire N881;
   wire N882;
   wire N883;
   wire N884;
   wire N885;
   wire N889;
   wire N945;
   wire N1110;
   wire N1111;
   wire N1112;
   wire N1113;
   wire N1114;
   wire N1489;
   wire N1490;
   wire N1781;
   wire N10025;
   wire N10101;
   wire N10102;
   wire N10103;
   wire N10104;
   wire N10109;
   wire N10110;
   wire N10111;
   wire N10112;
   wire N10350;
   wire N10351;
   wire N10352;
   wire N10353;
   wire N10574;
   wire N10575;
   wire N10576;
   wire N10628;
   wire N10632;
   wire N10641;
   wire N10704;
   wire N10706;
   wire N10711;
   wire N10712;
   wire N10713;
   wire N10714;
   wire N10715;
   wire N10716;
   wire N10717;
   wire N10718;
   wire N10729;
   wire N10759;
   wire N10760;
   wire N10761;
   wire N10762;
   wire N10763;
   wire N10827;
   wire N10837;
   wire N10838;
   wire N10839;
   wire N10840;
   wire N10868;
   wire N10869;
   wire N10870;
   wire N10871;
   wire N10905;
   wire N10906;
   wire N10907;
   wire N10908;
   wire N11333;
   wire N11334;
   wire N11340;
   wire N11342;
   wire N241_O;

   // map PI[] vector to DUT inputs and bidis
   assign N1 = PI[0];
   assign N5 = PI[1];
   assign N9 = PI[2];
   assign N12 = PI[3];
   assign N15 = PI[4];
   assign N18 = PI[5];
   assign N23 = PI[6];
   assign N26 = PI[7];
   assign N29 = PI[8];
   assign N32 = PI[9];
   assign N35 = PI[10];
   assign N38 = PI[11];
   assign N41 = PI[12];
   assign N44 = PI[13];
   assign N47 = PI[14];
   assign N50 = PI[15];
   assign N53 = PI[16];
   assign N54 = PI[17];
   assign N55 = PI[18];
   assign N56 = PI[19];
   assign N57 = PI[20];
   assign N58 = PI[21];
   assign N59 = PI[22];
   assign N60 = PI[23];
   assign N61 = PI[24];
   assign N62 = PI[25];
   assign N63 = PI[26];
   assign N64 = PI[27];
   assign N65 = PI[28];
   assign N66 = PI[29];
   assign N69 = PI[30];
   assign N70 = PI[31];
   assign N73 = PI[32];
   assign N74 = PI[33];
   assign N75 = PI[34];
   assign N76 = PI[35];
   assign N77 = PI[36];
   assign N78 = PI[37];
   assign N79 = PI[38];
   assign N80 = PI[39];
   assign N81 = PI[40];
   assign N82 = PI[41];
   assign N83 = PI[42];
   assign N84 = PI[43];
   assign N85 = PI[44];
   assign N86 = PI[45];
   assign N87 = PI[46];
   assign N88 = PI[47];
   assign N89 = PI[48];
   assign N94 = PI[49];
   assign N97 = PI[50];
   assign N100 = PI[51];
   assign N103 = PI[52];
   assign N106 = PI[53];
   assign N109 = PI[54];
   assign N110 = PI[55];
   assign N111 = PI[56];
   assign N112 = PI[57];
   assign N113 = PI[58];
   assign N114 = PI[59];
   assign N115 = PI[60];
   assign N118 = PI[61];
   assign N121 = PI[62];
   assign N124 = PI[63];
   assign N127 = PI[64];
   assign N130 = PI[65];
   assign N133 = PI[66];
   assign N134 = PI[67];
   assign N135 = PI[68];
   assign N138 = PI[69];
   assign N141 = PI[70];
   assign N144 = PI[71];
   assign N147 = PI[72];
   assign N150 = PI[73];
   assign N151 = PI[74];
   assign N152 = PI[75];
   assign N153 = PI[76];
   assign N154 = PI[77];
   assign N155 = PI[78];
   assign N156 = PI[79];
   assign N157 = PI[80];
   assign N158 = PI[81];
   assign N159 = PI[82];
   assign N160 = PI[83];
   assign N161 = PI[84];
   assign N162 = PI[85];
   assign N163 = PI[86];
   assign N164 = PI[87];
   assign N165 = PI[88];
   assign N166 = PI[89];
   assign N167 = PI[90];
   assign N168 = PI[91];
   assign N169 = PI[92];
   assign N170 = PI[93];
   assign N171 = PI[94];
   assign N172 = PI[95];
   assign N173 = PI[96];
   assign N174 = PI[97];
   assign N175 = PI[98];
   assign N176 = PI[99];
   assign N177 = PI[100];
   assign N178 = PI[101];
   assign N179 = PI[102];
   assign N180 = PI[103];
   assign N181 = PI[104];
   assign N182 = PI[105];
   assign N183 = PI[106];
   assign N184 = PI[107];
   assign N185 = PI[108];
   assign N186 = PI[109];
   assign N187 = PI[110];
   assign N188 = PI[111];
   assign N189 = PI[112];
   assign N190 = PI[113];
   assign N191 = PI[114];
   assign N192 = PI[115];
   assign N193 = PI[116];
   assign N194 = PI[117];
   assign N195 = PI[118];
   assign N196 = PI[119];
   assign N197 = PI[120];
   assign N198 = PI[121];
   assign N199 = PI[122];
   assign N200 = PI[123];
   assign N201 = PI[124];
   assign N202 = PI[125];
   assign N203 = PI[126];
   assign N204 = PI[127];
   assign N205 = PI[128];
   assign N206 = PI[129];
   assign N207 = PI[130];
   assign N208 = PI[131];
   assign N209 = PI[132];
   assign N210 = PI[133];
   assign N211 = PI[134];
   assign N212 = PI[135];
   assign N213 = PI[136];
   assign N214 = PI[137];
   assign N215 = PI[138];
   assign N216 = PI[139];
   assign N217 = PI[140];
   assign N218 = PI[141];
   assign N219 = PI[142];
   assign N220 = PI[143];
   assign N221 = PI[144];
   assign N222 = PI[145];
   assign N223 = PI[146];
   assign N224 = PI[147];
   assign N225 = PI[148];
   assign N226 = PI[149];
   assign N227 = PI[150];
   assign N228 = PI[151];
   assign N229 = PI[152];
   assign N230 = PI[153];
   assign N231 = PI[154];
   assign N232 = PI[155];
   assign N233 = PI[156];
   assign N234 = PI[157];
   assign N235 = PI[158];
   assign N236 = PI[159];
   assign N237 = PI[160];
   assign N238 = PI[161];
   assign N239 = PI[162];
   assign N240 = PI[163];
   assign N242 = PI[164];
   assign N245 = PI[165];
   assign N248 = PI[166];
   assign N251 = PI[167];
   assign N254 = PI[168];
   assign N257 = PI[169];
   assign N260 = PI[170];
   assign N263 = PI[171];
   assign N267 = PI[172];
   assign N271 = PI[173];
   assign N274 = PI[174];
   assign N277 = PI[175];
   assign N280 = PI[176];
   assign N283 = PI[177];
   assign N286 = PI[178];
   assign N289 = PI[179];
   assign N293 = PI[180];
   assign N296 = PI[181];
   assign N299 = PI[182];
   assign N303 = PI[183];
   assign N307 = PI[184];
   assign N310 = PI[185];
   assign N313 = PI[186];
   assign N316 = PI[187];
   assign N319 = PI[188];
   assign N322 = PI[189];
   assign N325 = PI[190];
   assign N328 = PI[191];
   assign N331 = PI[192];
   assign N334 = PI[193];
   assign N337 = PI[194];
   assign N340 = PI[195];
   assign N343 = PI[196];
   assign N346 = PI[197];
   assign N349 = PI[198];
   assign N352 = PI[199];
   assign N355 = PI[200];
   assign N358 = PI[201];
   assign N361 = PI[202];
   assign N364 = PI[203];
   assign N367 = PI[204];
   assign N382 = PI[205];
   assign N241_I = PI[206];

   // map DUT outputs and bidis to PO[] vector
   assign
      PO[0] = N387 ,
      PO[1] = N388 ,
      PO[2] = N478 ,
      PO[3] = N482 ,
      PO[4] = N484 ,
      PO[5] = N486 ,
      PO[6] = N489 ,
      PO[7] = N492 ,
      PO[8] = N501 ,
      PO[9] = N505 ,
      PO[10] = N507 ,
      PO[11] = N509 ,
      PO[12] = N511 ,
      PO[13] = N513 ,
      PO[14] = N515 ,
      PO[15] = N517 ,
      PO[16] = N519 ,
      PO[17] = N535 ,
      PO[18] = N537 ,
      PO[19] = N539 ,
      PO[20] = N541 ,
      PO[21] = N543 ,
      PO[22] = N545 ,
      PO[23] = N547 ,
      PO[24] = N549 ,
      PO[25] = N551 ,
      PO[26] = N553 ,
      PO[27] = N556 ,
      PO[28] = N559 ,
      PO[29] = N561 ,
      PO[30] = N563 ,
      PO[31] = N565 ;
   assign
      PO[32] = N567 ,
      PO[33] = N569 ,
      PO[34] = N571 ,
      PO[35] = N573 ,
      PO[36] = N582 ,
      PO[37] = N643 ,
      PO[38] = N707 ,
      PO[39] = N813 ,
      PO[40] = N881 ,
      PO[41] = N882 ,
      PO[42] = N883 ,
      PO[43] = N884 ,
      PO[44] = N885 ,
      PO[45] = N889 ,
      PO[46] = N945 ,
      PO[47] = N1110 ,
      PO[48] = N1111 ,
      PO[49] = N1112 ,
      PO[50] = N1113 ,
      PO[51] = N1114 ,
      PO[52] = N1489 ,
      PO[53] = N1490 ,
      PO[54] = N1781 ,
      PO[55] = N10025 ,
      PO[56] = N10101 ,
      PO[57] = N10102 ,
      PO[58] = N10103 ,
      PO[59] = N10104 ,
      PO[60] = N10109 ,
      PO[61] = N10110 ,
      PO[62] = N10111 ,
      PO[63] = N10112 ;
   assign
      PO[64] = N10350 ,
      PO[65] = N10351 ,
      PO[66] = N10352 ,
      PO[67] = N10353 ,
      PO[68] = N10574 ,
      PO[69] = N10575 ,
      PO[70] = N10576 ,
      PO[71] = N10628 ,
      PO[72] = N10632 ,
      PO[73] = N10641 ,
      PO[74] = N10704 ,
      PO[75] = N10706 ,
      PO[76] = N10711 ,
      PO[77] = N10712 ,
      PO[78] = N10713 ,
      PO[79] = N10714 ,
      PO[80] = N10715 ,
      PO[81] = N10716 ,
      PO[82] = N10717 ,
      PO[83] = N10718 ,
      PO[84] = N10729 ,
      PO[85] = N10759 ,
      PO[86] = N10760 ,
      PO[87] = N10761 ,
      PO[88] = N10762 ,
      PO[89] = N10763 ,
      PO[90] = N10827 ,
      PO[91] = N10837 ,
      PO[92] = N10838 ,
      PO[93] = N10839 ,
      PO[94] = N10840 ,
      PO[95] = N10868 ;
   assign
      PO[96] = N10869 ,
      PO[97] = N10870 ,
      PO[98] = N10871 ,
      PO[99] = N10905 ,
      PO[100] = N10906 ,
      PO[101] = N10907 ,
      PO[102] = N10908 ,
      PO[103] = N11333 ,
      PO[104] = N11334 ,
      PO[105] = N11340 ,
      PO[106] = N11342 ,
      PO[107] = N241_O ;

   // instantiate the design into the testbench
   c7552 dut (
      .N1(N1),
      .N5(N5),
      .N9(N9),
      .N12(N12),
      .N15(N15),
      .N18(N18),
      .N23(N23),
      .N26(N26),
      .N29(N29),
      .N32(N32),
      .N35(N35),
      .N38(N38),
      .N41(N41),
      .N44(N44),
      .N47(N47),
      .N50(N50),
      .N53(N53),
      .N54(N54),
      .N55(N55),
      .N56(N56),
      .N57(N57),
      .N58(N58),
      .N59(N59),
      .N60(N60),
      .N61(N61),
      .N62(N62),
      .N63(N63),
      .N64(N64),
      .N65(N65),
      .N66(N66),
      .N69(N69),
      .N70(N70),
      .N73(N73),
      .N74(N74),
      .N75(N75),
      .N76(N76),
      .N77(N77),
      .N78(N78),
      .N79(N79),
      .N80(N80),
      .N81(N81),
      .N82(N82),
      .N83(N83),
      .N84(N84),
      .N85(N85),
      .N86(N86),
      .N87(N87),
      .N88(N88),
      .N89(N89),
      .N94(N94),
      .N97(N97),
      .N100(N100),
      .N103(N103),
      .N106(N106),
      .N109(N109),
      .N110(N110),
      .N111(N111),
      .N112(N112),
      .N113(N113),
      .N114(N114),
      .N115(N115),
      .N118(N118),
      .N121(N121),
      .N124(N124),
      .N127(N127),
      .N130(N130),
      .N133(N133),
      .N134(N134),
      .N135(N135),
      .N138(N138),
      .N141(N141),
      .N144(N144),
      .N147(N147),
      .N150(N150),
      .N151(N151),
      .N152(N152),
      .N153(N153),
      .N154(N154),
      .N155(N155),
      .N156(N156),
      .N157(N157),
      .N158(N158),
      .N159(N159),
      .N160(N160),
      .N161(N161),
      .N162(N162),
      .N163(N163),
      .N164(N164),
      .N165(N165),
      .N166(N166),
      .N167(N167),
      .N168(N168),
      .N169(N169),
      .N170(N170),
      .N171(N171),
      .N172(N172),
      .N173(N173),
      .N174(N174),
      .N175(N175),
      .N176(N176),
      .N177(N177),
      .N178(N178),
      .N179(N179),
      .N180(N180),
      .N181(N181),
      .N182(N182),
      .N183(N183),
      .N184(N184),
      .N185(N185),
      .N186(N186),
      .N187(N187),
      .N188(N188),
      .N189(N189),
      .N190(N190),
      .N191(N191),
      .N192(N192),
      .N193(N193),
      .N194(N194),
      .N195(N195),
      .N196(N196),
      .N197(N197),
      .N198(N198),
      .N199(N199),
      .N200(N200),
      .N201(N201),
      .N202(N202),
      .N203(N203),
      .N204(N204),
      .N205(N205),
      .N206(N206),
      .N207(N207),
      .N208(N208),
      .N209(N209),
      .N210(N210),
      .N211(N211),
      .N212(N212),
      .N213(N213),
      .N214(N214),
      .N215(N215),
      .N216(N216),
      .N217(N217),
      .N218(N218),
      .N219(N219),
      .N220(N220),
      .N221(N221),
      .N222(N222),
      .N223(N223),
      .N224(N224),
      .N225(N225),
      .N226(N226),
      .N227(N227),
      .N228(N228),
      .N229(N229),
      .N230(N230),
      .N231(N231),
      .N232(N232),
      .N233(N233),
      .N234(N234),
      .N235(N235),
      .N236(N236),
      .N237(N237),
      .N238(N238),
      .N239(N239),
      .N240(N240),
      .N242(N242),
      .N245(N245),
      .N248(N248),
      .N251(N251),
      .N254(N254),
      .N257(N257),
      .N260(N260),
      .N263(N263),
      .N267(N267),
      .N271(N271),
      .N274(N274),
      .N277(N277),
      .N280(N280),
      .N283(N283),
      .N286(N286),
      .N289(N289),
      .N293(N293),
      .N296(N296),
      .N299(N299),
      .N303(N303),
      .N307(N307),
      .N310(N310),
      .N313(N313),
      .N316(N316),
      .N319(N319),
      .N322(N322),
      .N325(N325),
      .N328(N328),
      .N331(N331),
      .N334(N334),
      .N337(N337),
      .N340(N340),
      .N343(N343),
      .N346(N346),
      .N349(N349),
      .N352(N352),
      .N355(N355),
      .N358(N358),
      .N361(N361),
      .N364(N364),
      .N367(N367),
      .N382(N382),
      .N241_I(N241_I),
      .N387(N387),
      .N388(N388),
      .N478(N478),
      .N482(N482),
      .N484(N484),
      .N486(N486),
      .N489(N489),
      .N492(N492),
      .N501(N501),
      .N505(N505),
      .N507(N507),
      .N509(N509),
      .N511(N511),
      .N513(N513),
      .N515(N515),
      .N517(N517),
      .N519(N519),
      .N535(N535),
      .N537(N537),
      .N539(N539),
      .N541(N541),
      .N543(N543),
      .N545(N545),
      .N547(N547),
      .N549(N549),
      .N551(N551),
      .N553(N553),
      .N556(N556),
      .N559(N559),
      .N561(N561),
      .N563(N563),
      .N565(N565),
      .N567(N567),
      .N569(N569),
      .N571(N571),
      .N573(N573),
      .N582(N582),
      .N643(N643),
      .N707(N707),
      .N813(N813),
      .N881(N881),
      .N882(N882),
      .N883(N883),
      .N884(N884),
      .N885(N885),
      .N889(N889),
      .N945(N945),
      .N1110(N1110),
      .N1111(N1111),
      .N1112(N1112),
      .N1113(N1113),
      .N1114(N1114),
      .N1489(N1489),
      .N1490(N1490),
      .N1781(N1781),
      .N10025(N10025),
      .N10101(N10101),
      .N10102(N10102),
      .N10103(N10103),
      .N10104(N10104),
      .N10109(N10109),
      .N10110(N10110),
      .N10111(N10111),
      .N10112(N10112),
      .N10350(N10350),
      .N10351(N10351),
      .N10352(N10352),
      .N10353(N10353),
      .N10574(N10574),
      .N10575(N10575),
      .N10576(N10576),
      .N10628(N10628),
      .N10632(N10632),
      .N10641(N10641),
      .N10704(N10704),
      .N10706(N10706),
      .N10711(N10711),
      .N10712(N10712),
      .N10713(N10713),
      .N10714(N10714),
      .N10715(N10715),
      .N10716(N10716),
      .N10717(N10717),
      .N10718(N10718),
      .N10729(N10729),
      .N10759(N10759),
      .N10760(N10760),
      .N10761(N10761),
      .N10762(N10762),
      .N10763(N10763),
      .N10827(N10827),
      .N10837(N10837),
      .N10838(N10838),
      .N10839(N10839),
      .N10840(N10840),
      .N10868(N10868),
      .N10869(N10869),
      .N10870(N10870),
      .N10871(N10871),
      .N10905(N10905),
      .N10906(N10906),
      .N10907(N10907),
      .N10908(N10908),
      .N11333(N11333),
      .N11334(N11334),
      .N11340(N11340),
      .N11342(N11342),
      .N241_O(N241_O)   );


   integer errshown;
   event measurePO;
   always @ measurePO begin
      if (((XPCT&MASK) !== (ALLPOS&MASK)) || (XPCT !== (~(~XPCT)))) begin
         errshown = 0;
         for (bit = 0; bit < NOUTPUTS; bit=bit + 1) begin
            if (MASK[bit]==1'b1) begin
               if (XPCT[bit] !== ALLPOS[bit]) begin
                  if (errshown==0) $display("\n// *** ERROR during capture pattern %0d, T=%t", pattern, $time);
                  $display("  %0d %0s (exp=%b, got=%b)", pattern, POnames[bit], XPCT[bit], ALLPOS[bit]);
                  nofails = nofails + 1; errshown = 1;
               end
            end
         end
      end
   end

   event forcePI_default_WFT;
   always @ forcePI_default_WFT begin
      PI = ALLPIS;
   end
   event measurePO_default_WFT;
   always @ measurePO_default_WFT begin
      #40;
      ALLPOS = PO;
      #0; #0 -> measurePO;
      `ifdef tmax_iddq
         #0; ->IDDQ;
      `endif
   end

   always @ IDDQ begin
   `ifdef tmax_iddq
      $ssi_iddq("strobe_try");
      $ssi_iddq("status drivers leaky AAA_tmax_testbench_1_16.leaky");
   `endif
   end

   event capture;
   always @ capture begin
      ->forcePI_default_WFT;
      #100; ->measurePO_default_WFT;
   end


   initial begin

      //
      // --- establish a default time format for %t
      //
      $timeformat(-9,2," ns",18);

      //
      // --- default verbosity to 2 but also allow user override by
      //     using '+define+tmax_msg=N' on verilog compile line.
      //
      `ifdef tmax_msg
         verbose = `tmax_msg ;
      `else
         verbose = 2 ;
      `endif

      //
      // --- default pattern reporting interval to 5 but also allow user
      //     override by using '+define+tmax_rpt=N' on verilog compile line.
      //
      `ifdef tmax_rpt
         report_interval = `tmax_rpt ;
      `else
         report_interval = 5 ;
      `endif

      //
      // --- support generating Extened VCD output by using
      //     '+define+tmax_vcde' on verilog compile line.
      //
      `ifdef tmax_vcde
         // extended VCD, see IEEE Verilog P1364.1-1999 Draft 2
         if (verbose >= 2) $display("// %t : opening Extended VCD output file", $time);
         $dumpports( dut, "sim_vcde.out");
      `endif

      //
      // --- IDDQ PLI initialization
      //     User may activite by using '+define+tmax_iddq' on verilog compile line.
      //     Or by defining `tmax_iddq in this file.
      //
      `ifdef tmax_iddq
         if (verbose >= 3) $display("// %t : Initializing IDDQ PLI", $time);
         $ssi_iddq("dut AAA_tmax_testbench_1_16.dut");
         $ssi_iddq("verb on");
         $ssi_iddq("cycle 0");
         //
         // --- User may select one of the following two methods for fault seeding:
         //     #1 faults seeded by PLI (default)
         //     #2 faults supplied in a file
         //     Comment out the unused lines as needed (precede with '//').
         //     Replace the 'FAULTLIST_FILE' string with the actual file pathname.
         //
         $ssi_iddq("seed SA AAA_tmax_testbench_1_16.dut");   // no file, faults seeded by PLI
         //
         // $ssi_iddq("scope AAA_tmax_testbench_1_16.dut");   // set scope for faults from a file
         // $ssi_iddq("read_tmax FAULTLIST_FILE"); // read faults from a file
         //
      `endif

      POnames[0] = "N387";
      POnames[1] = "N388";
      POnames[2] = "N478";
      POnames[3] = "N482";
      POnames[4] = "N484";
      POnames[5] = "N486";
      POnames[6] = "N489";
      POnames[7] = "N492";
      POnames[8] = "N501";
      POnames[9] = "N505";
      POnames[10] = "N507";
      POnames[11] = "N509";
      POnames[12] = "N511";
      POnames[13] = "N513";
      POnames[14] = "N515";
      POnames[15] = "N517";
      POnames[16] = "N519";
      POnames[17] = "N535";
      POnames[18] = "N537";
      POnames[19] = "N539";
      POnames[20] = "N541";
      POnames[21] = "N543";
      POnames[22] = "N545";
      POnames[23] = "N547";
      POnames[24] = "N549";
      POnames[25] = "N551";
      POnames[26] = "N553";
      POnames[27] = "N556";
      POnames[28] = "N559";
      POnames[29] = "N561";
      POnames[30] = "N563";
      POnames[31] = "N565";
      POnames[32] = "N567";
      POnames[33] = "N569";
      POnames[34] = "N571";
      POnames[35] = "N573";
      POnames[36] = "N582";
      POnames[37] = "N643";
      POnames[38] = "N707";
      POnames[39] = "N813";
      POnames[40] = "N881";
      POnames[41] = "N882";
      POnames[42] = "N883";
      POnames[43] = "N884";
      POnames[44] = "N885";
      POnames[45] = "N889";
      POnames[46] = "N945";
      POnames[47] = "N1110";
      POnames[48] = "N1111";
      POnames[49] = "N1112";
      POnames[50] = "N1113";
      POnames[51] = "N1114";
      POnames[52] = "N1489";
      POnames[53] = "N1490";
      POnames[54] = "N1781";
      POnames[55] = "N10025";
      POnames[56] = "N10101";
      POnames[57] = "N10102";
      POnames[58] = "N10103";
      POnames[59] = "N10104";
      POnames[60] = "N10109";
      POnames[61] = "N10110";
      POnames[62] = "N10111";
      POnames[63] = "N10112";
      POnames[64] = "N10350";
      POnames[65] = "N10351";
      POnames[66] = "N10352";
      POnames[67] = "N10353";
      POnames[68] = "N10574";
      POnames[69] = "N10575";
      POnames[70] = "N10576";
      POnames[71] = "N10628";
      POnames[72] = "N10632";
      POnames[73] = "N10641";
      POnames[74] = "N10704";
      POnames[75] = "N10706";
      POnames[76] = "N10711";
      POnames[77] = "N10712";
      POnames[78] = "N10713";
      POnames[79] = "N10714";
      POnames[80] = "N10715";
      POnames[81] = "N10716";
      POnames[82] = "N10717";
      POnames[83] = "N10718";
      POnames[84] = "N10729";
      POnames[85] = "N10759";
      POnames[86] = "N10760";
      POnames[87] = "N10761";
      POnames[88] = "N10762";
      POnames[89] = "N10763";
      POnames[90] = "N10827";
      POnames[91] = "N10837";
      POnames[92] = "N10838";
      POnames[93] = "N10839";
      POnames[94] = "N10840";
      POnames[95] = "N10868";
      POnames[96] = "N10869";
      POnames[97] = "N10870";
      POnames[98] = "N10871";
      POnames[99] = "N10905";
      POnames[100] = "N10906";
      POnames[101] = "N10907";
      POnames[102] = "N10908";
      POnames[103] = "N11333";
      POnames[104] = "N11334";
      POnames[105] = "N11340";
      POnames[106] = "N11342";
      POnames[107] = "N241_O";
      nofails = 0; pattern = -1; lastpattern = 0;
      prev_pat = -2; error_banner = -2;
      /*** No test setup procedure ***/


      /*** Non-scan test ***/

      if (verbose >= 1) $display("// %t : Begin patterns, first pattern = 0", $time);
pattern = 0; // 0
ALLPIS = 207'b111000001101100000110111100011011101001101000110101101001100011001100010111001001110001011010000101111101110000111100100101110001110011100100000001011010111110100011110101001111110011110111111011000011001100;
XPCT = 108'b111101001111001111011111101100011001101011111111111111111111001011011111011100010100110001011111101000011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 200

pattern = 1; // 200
ALLPIS = 207'b111100000110110000011011110001101110100110100011010110100110001100110001011100100111000101101000010111110111000011110010010111000111001110010000000101101011111010001111010100111111001111011111101100001100110;
XPCT = 108'b111010101111100111101111110100001100111111111101111111000000101001000100101000101011100011111000101100011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 400

pattern = 2; // 400
ALLPIS = 207'b100110001110111000111010011011101010011110010111000110011111011111111010010111011101101001100100100100010101100110011101100101101101111011101000001001100010001001011001000011100001111001010000101110011111111;
XPCT = 108'b110000011000111100101000010110011111010111111100000001100000011110111110101000111111101000011000011110010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 600

pattern = 3; // 600
ALLPIS = 207'b001011001010111100101010101110101000000010001101001110000011110110011111110010100000111111100010111101100100110100101010011100111000100001010100001111100110110000110010001000001110100010010111001111010110011;
XPCT = 108'b001001000111010001001011100111010110000111111001011010010000010101111110110010001101101000111110011101001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 800

pattern = 4; // 800
ALLPIS = 207'b011101101000111110100010110100001001001100000000001010001101100010101101000000011110010100100001110001011100011101110001100000010010001100001010001100100100101100000111101101111001001111110100111111110010101;
XPCT = 108'b001101101100100111111010011111110010111111111001111110000000000101101110101011000110100011111111100001101001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1000

pattern = 5; // 1000
ALLPIS = 207'b001110110100011111010001011010000100100110000000000101000110110001010110100000001111001010010000111000101110001110111000110000001001000110000101000110010010010110000011110110111100100111111010011111111001010;
XPCT = 108'b001110111110010011111101001111111001011101111011011010000000111011110100101011011000100110100001000110010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1200

pattern = 6; // 1200
ALLPIS = 207'b111111010111101111011111001110011111011110000110101111101111000001001001101001001001101110011000110011111001000000111000110110001010111111100010101000011110111111011111010010100000001101000010010111100101001;
XPCT = 108'b111010011000000110100001001011100101010111111111011011111111111000101111100100011001110100111000000000000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1400

pattern = 7; // 1400
ALLPIS = 207'b011111101011110111101111100111001111101111000011010111110111100000100100110100100100110111001100011001111100100000011100011011000101011111110001010100001111011111101111101001010000000110100001001011110010100;
XPCT = 108'b001101000000000011010000100111110010011011111011011010001111111010111111100100110100111000011000101000011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1600

pattern = 8; // 1600
ALLPIS = 207'b010111111000011011000000010000111010111010100111000110110111101001110000100011011100010000110110100011010000010111101010100011101100110011011000100001010000011011101001011101010110011101101111111101100000110;
XPCT = 108'b000011100011001110110111111101100000011111111001011010000000111000011110111001010000101111111111010000100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 1800

pattern = 9; // 1800
ALLPIS = 207'b001011111100001101100000001000011101011101010011100011011011110100111000010001101110001000011011010001101000001011110101010001110110011001101100010000101000001101110100101110101011001110110111111110110000011;
XPCT = 108'b000101111101100111011011111110110000000101111011010000010000000100010110011000011010101010100000010000000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2000

pattern = 10; // 2000
ALLPIS = 207'b100101111110000110110000000100001110101110101001110001101101111010011100001000110111000100001101101000110100000101111010101000111011001100110110001000010100000110111010010111010101100111011011111111011000001;
XPCT = 108'b111010110010110011101101111111011000101101111110101111010000111100001110011011011100101001011111100011000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2200

pattern = 11; // 2200
ALLPIS = 207'b001010110010100011101111100001011010011010010010010101111010100100101100111101010101101001010110011011110100000101011001111010010011111010111011001111011101110111000011100010010100101101010010100111110101100;
XPCT = 108'b001100010010010110101001010011110101011111111011011010001111010001111111101110101100110010100000010111011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2400

pattern = 12; // 2400
ALLPIS = 207'b111101010100110001000000010011110000000000001111100111110001001011110100100111100100111111111011100010010100000101001000010011000111100001111101101100111001001111111111011000110100001000010110001011100011010;
XPCT = 108'b111011001010000100001011000111100011111011111111111111110000010000111110000000010001101100111110101101000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2600

pattern = 13; // 2600
ALLPIS = 207'b011110101010011000100000001001111000000000000111110011111000100101111010010011110010011111111101110001001010000010100100001001100011110000111110110110011100100111111111101100011010000100001011000101110001101;
XPCT = 108'b001101100101000010000101100001110001011111111011011010000000100100101110100011100100100111111111011000000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 2800

pattern = 14; // 2800
ALLPIS = 207'b110111011000101100100111100111100001001101000101010100110000001011011111110000110111000100101110010111001011000110110110101010111111100100111111010000011001100111100001011111110011011100111010111010100001010;
XPCT = 108'b110011111001101110011101011110100001011011111101011011010000111110001110111010100110100100000001011010010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3000

pattern = 15; // 3000
ALLPIS = 207'b111011101100010110010011110011110000100110100010101010011000000101101111111000011011100010010111001011100101100011011011010101011111110010011111101000001100110011110000101111111001101110011101011101010000101;
XPCT = 108'b110101111100110111001110101101010000001111111101011011001001010110001110001100100000110100100001101110111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3200

pattern = 16; // 3200
ALLPIS = 207'b100101111011101011111110011010100101011110010111111000000000011011010101000101000011111010011011001010011100110110001001000100100001100101101111111111010001101101100110111110000010101001110001110110110001110;
XPCT = 108'b111111110001010100111000111010110001100111111101111111100110101010001101000011111001101110111110001011101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3400

pattern = 17; // 3400
ALLPIS = 207'b001010110000010101001000101110001111100010001101010001001100010100001000011011101111110110011101001010100000011100100000001100011110101110010111110100111111000010101101110110111111001010000111100011000001011;
XPCT = 108'b000110111111100101000011110011000001011011110010001010010000110111001110000011001000101010000111111101111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3600

pattern = 18; // 3600
ALLPIS = 207'b100101011000001010100100010111000111110001000110101000100110001010000100001101110111111011001110100101010000001110010000000110001111010111001011111010011111100001010110111011011111100101000011110001100000101;
XPCT = 108'b111111010111110010100001111001100000101001111101111111100000000111111110011010001110101101011110100111111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 3800

pattern = 19; // 3800
ALLPIS = 207'b110010101100000101010010001011100011111000100011010100010011000101000010000110111011111101100111010010101000000111001000000011000111101011100101111101001111110000101011011101101111110010100001111000110000010;
XPCT = 108'b111011101111111001010000111100110000010011111101011011110000001111111110000010010011101011111110101110101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4000

pattern = 20; // 4000
ALLPIS = 207'b111001010110000010101001000101110001111100010001101010001001100010100001000011011101111110110011101001010100000011100100000001100011110101110010111110100111111000010101101110110111111001010000111100011000001;
XPCT = 108'b110101111011111100101000011100011000111111111101111111110000010100110110101011101110100101111110101101010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4200

pattern = 21; // 4200
ALLPIS = 207'b111100101011000001010100100010111000111110001000110101000100110001010000100001101110111111011001110100101010000001110010000000110001111010111001011111010011111100001010110111011011111100101000011110001100000;
XPCT = 108'b111110110101111110010100001110001100101111111111111111111111111100001111110100101000110000011000001111010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4400

pattern = 22; // 4400
ALLPIS = 207'b000110011000000000011101110010000001010010000010110111101110000001001010101001111001010100111100010101111011000111011101101110010110100001111100100100111110001010011011110010010011100000101011010111011111100;
XPCT = 108'b001110010001110000010101101011011111011111111010001010001111011011101111100111111000111101000000110000010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4600

pattern = 23; // 4600
ALLPIS = 207'b011011000001100000111001011010011101100100000111110110111011011001000111101101110010100001001110100101010011100100001010011001000101001100011110011001001000110001010011010000110111101110101010110011110110010;
XPCT = 108'b001010001011110111010101011011110110011011111001011010011111101101011111000101001100111001011001010001000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 4800

pattern = 24; // 4800
ALLPIS = 207'b010101101101010000101011001110010011111111000101010110010001110101000001001111110111011011110111111101000111110101100001100010101100111010101111000111110011101100110111000001100101101001101010000001100010101;
XPCT = 108'b001000001010110100110101000001100010110011101001111110001111011111011111101111011010111001111110001100011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5000

pattern = 25; // 5000
ALLPIS = 207'b101010110110101000010101100111001001111111100010101011001000111010100000100111111011101101111011111110100011111010110000110001010110011101010111100011111001110110011011100000110010110100110101000000110001010;
XPCT = 108'b111100001001011010011010100000110001011001111110001011101001001100001110001101001100110100100000001001111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5200

pattern = 26; // 5200
ALLPIS = 207'b101101010110110100111101010000111001110010110111111000101000000100110010101010110011111101101101010000111111111010111100110110100101010010001011111010101011001111010011011001100111000100100101111000000001001;
XPCT = 108'b111011001011100010010010111100000001110011101101110101110000010111101110101001010011100111011111010011111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5400

pattern = 27; // 5400
ALLPIS = 207'b110110101011011010011110101000011100111001011011111100010100000010011001010101011001111110110110101000011111111101011110011011010010101001000101111101010101100111101001101100110011100010010010111100000000100;
XPCT = 108'b110101101001110001001001011100000000011111101101011011101111001111011111100100010110111110011111010000101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5600

pattern = 28; // 5600
ALLPIS = 207'b000011011000001101111000110111010011010001101011010011000110011000101110010011100010110100001011111011100001111001001011100011100111001000000010110101111101000111101010011111100111101111110110000110011001110;
XPCT = 108'b001011111011110111111011000010011001000111111010001010000000110000101110000001000010100000100001011000100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 5800

pattern = 29; // 5800
ALLPIS = 207'b000001101100000110111100011011101001101000110101101001100011001100010111001001110001011010000101111101110000111100100101110001110011100100000001011010111110100011110101001111110011110111111011000011001100111;
XPCT = 108'b000001111001111011111101100011001100111011111011111110000000110001101110010001010101101011000000111001000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6000

pattern = 30; // 6000
ALLPIS = 207'b100000110110000011011110001101110100110100011010110100110001100110001011100100111000101101000010111110111000011110010010111000111001110010000000101101011111010001111010100111111001111011111101100001100110011;
XPCT = 108'b111100111100111101111110110001100110101011111100101111100000011001110100010001011110101000000111100010000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6200

pattern = 31; // 6200
ALLPIS = 207'b110000011011000001101111000110111010011010001101011010011000110011000101110010011100010110100001011111011100001111001001011100011100111001000000010110101111101000111101010011111100111101111110110000110011001;
XPCT = 108'b110010011110011110111111011000110011111011110101111111001111101101011111100101111011110000011110111010010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6400

pattern = 32; // 6400
ALLPIS = 207'b111010001001101010011110001011001000100000010110011000110001000110010000110011010010110101001001001010011101111000001000001111100100110110100111011111110010100101010111111001000010010010100010101010001110000;
XPCT = 108'b111111000001001001010001010110001110010010111101011011001111000000011111100101000010111101011111010000100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6600

pattern = 33; // 6600
ALLPIS = 207'b110100101011110000111001101001111010101000010011111110111101010111110100111111100110011000011011011000111010100110001010001100011101111011001110101000001110001100000010000111010010110110001010000000101101100;
XPCT = 108'b111000110001011011000101000000101101101011010101111111111111100111100101111101001111110100111111111110100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 6800

pattern = 34; // 6800
ALLPIS = 207'b000000011100010010000010111111110101110100011111100111101111101101101010101100100001111001000100100110000000101011001101001001101010001011000000001011110101100011010110111010101011001001100111101010011000110;
XPCT = 108'b001111011101100100110011110110011000100001111011111110010000000101101110111011110000101010011001011100001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7000

pattern = 35; // 7000
ALLPIS = 207'b011010000111100011011111010100110010011010011001101011000110110000100101100101000010001001101011011001011101101101101110101011010001110011000111011010001000010100111100100100010111110110010001011111000010011;
XPCT = 108'b000100100011111011001000101111000010001111111011011010001111011001101111110111001100110011111001101111001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7200

pattern = 36; // 7200
ALLPIS = 207'b101100101000010010101001111110000100000110110000000010000000101010011001101010000010010111010011111100001010100011010011100101010000101010010110101001010000100000011000110000000111101111000110111101111110100;
XPCT = 108'b110110000011110111100011011101111110100111111100101111010000010001011110010010001010100010011110101100010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7400

pattern = 37; // 7400
ALLPIS = 207'b110110010100001001010100111111000010000011011000000001000000010101001100110101000001001011101001111110000101010001101001110010101000010101001011010100101000010000001100011000000011110111100011011110111111010;
XPCT = 108'b110011000001111011110001101110111111000111111111011011101001000010101110011100010001110100100001010101011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7600

pattern = 38; // 7600
ALLPIS = 207'b100001000011101110110100010100101001100001111010011000010001001100110110101001110010010000111101110101011111010000111100110110110000111100000010110101100110101101010001110101000011101001010011000101010001101;
XPCT = 108'b110110100001110100101001100001010001110101111101110101001111101101111111100101101011110001111001010001011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 7800

pattern = 39; // 7800
ALLPIS = 207'b010000100001110111011010001010010100110000111101001100001000100110011011010100111001001000011110111010101111101000011110011011011000011110000001011010110011010110101000111010100001110100101001100010101000110;
XPCT = 108'b000111011000111010010100110010101000100011111001111110011111111101111111010101100010110100000111100001000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8000

pattern = 40; // 8000
ALLPIS = 207'b101000010000111011101101000101001010011000011110100110000100010011001101101010011100100100001111011101010111110100001111001101101100001111000000101101011001101011010100011101010000111010010100110001010100011;
XPCT = 108'b110011100000011101001010011001010100101011101101111111000110000011110101010011110011101000011111110010100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8200

pattern = 41; // 8200
ALLPIS = 207'b001110000001110111101000101001101101101100011001001011110011001111110110000110011100100111001110100100110110000010001111101001010010110001000111001001011110010000111101110111101010001111101000110010100100001;
XPCT = 108'b000110111101000111110100011010100100010011011010000000011111001010111111001111001000110011111001111100111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8400

pattern = 42; // 8400
ALLPIS = 207'b111101001001010001101010011111111110010110011010111101001000100001101011110000011100100110101110011000000110111001001111111011001101101110000100111011011101101101001001000010110111010101010110110011011100000;
XPCT = 108'b110000011011101010101011011011011100111011101111111111011111001010011111001101011101110101111001111111111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8600

pattern = 43; // 8600
ALLPIS = 207'b011110100100101000110101001111111111001011001101011110100100010000110101111000001110010011010111001100000011011100100111111101100110110111000010011101101110110110100100100001011011101010101011011001101110000;
XPCT = 108'b000100000101110101010101101101101110001011110001011010000000011111011110010001101110101010011110101001111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 8800

pattern = 44; // 8800
ALLPIS = 207'b010101011011111110000100101100110111000101110000110111100011001110001010001111010101111100100010101100011100010110011011110001010111101101000110010001000101111110000101101001101111100111110111000110111001000;
XPCT = 108'b000101001111110011111011100010111001110111111011111110011111001001001111000101101001110011111000011111110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9000

pattern = 45; // 9000
ALLPIS = 207'b001010101101111111000010010110011011100010111000011011110001100111000101000111101010111110010001010110001110001011001101111000101011110110100011001000100010111111000010110100110111110011111011100011011100100;
XPCT = 108'b001110101011111001111101110011011100001001111011011010001111011000001111110111001000111011011110000001111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9200

pattern = 46; // 9200
ALLPIS = 207'b011111011111010101111111000000000101010001001010010101001001110101110010010000100111101010000001100001011010111101101110110011110001001101110110111011100011111010110110100011011001101011011111011011100000010;
XPCT = 108'b001100010100110101101111101111100000001011111011011010011111101100111111111111011100111010000000100101110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9400

pattern = 47; // 9400
ALLPIS = 207'b110101100110000000100001101011001010001000110011010010010101111100101001111011000001000000001001111010110000100110111111010110011100010000011100000010000011011000001100101000101110100111001101000111111110001;
XPCT = 108'b110101001111010011100110100011111110100111111101111111010000101110101110001010101000100010011110011100000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9600

pattern = 48; // 9600
ALLPIS = 207'b111010110011000000010000110101100101000100011001101001001010111110010100111101100000100000000100111101011000010011011111101011001110001000001110000001000001101100000110010100010111010011100110100011111111000;
XPCT = 108'b111010100011101001110011010011111111001011111111011011001111110000001111111110101001111100111110110100100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 9800

pattern = 49; // 9800
ALLPIS = 207'b111101011001100000001000011010110010100010001100110100100101011111001010011110110000010000000010011110101100001001101111110101100111000100000111000000100000110110000011001010001011101001110011010001111111100;
XPCT = 108'b111001010101110100111001101001111111110011111101111111001111001110001111000100110111111010111000001110011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10000

pattern = 50; // 10000
ALLPIS = 207'b011110101100110000000100001101011001010001000110011010010010101111100101001111011000001000000001001111010110000100110111111010110011100010000011100000010000011011000001100101000101110100111001101000111111110;
XPCT = 108'b000100100010111010011100110100111111010011111001011010010000011000011110100010001110100100011001011101001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10200

pattern = 51; // 10200
ALLPIS = 207'b101111010110011000000010000110101100101000100011001101001001010111110010100111101100000100000000100111101011000010011011111101011001110001000001110000001000001101100000110010100010111010011100110100011111111;
XPCT = 108'b110110011001011101001110011000011111000101111111010001000000111100110110110011111000101000000110111011110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10400

pattern = 52; // 10400
ALLPIS = 207'b101101100010100110011111001000011110110100000111111110010101101101101001100000100100110111001001011001101000011001000101110001001000001110000111100111110110100011100111100000010011001111101100110000000001111;
XPCT = 108'b111100000001100111110110011000000001111011111101111111000000011011011000100001111110100011111110110011010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10600

pattern = 53; // 10600
ALLPIS = 207'b101100111000111001010001101111000111111010010101100111111011110000100100000011000000101110101101100110101001110100101010110111000000110001100100101100001001110100100100001001001011110101010100110010001110111;
XPCT = 108'b110001000101111010101010011010001110100001111111111111100000010111001110010001000101100100011110111000110111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 10800

pattern = 54; // 10800
ALLPIS = 207'b110110001010111011011011011110010101101110101110010101100110011111000001011001011001010001001111111100100100100001001110101010000010010111001010100100111011001111100010111110110011110100000100011001100100101;
XPCT = 108'b111111111001111010000010001101100100001011111111011011011111100101101111010111010000110011100001000111100101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11000

pattern = 55; // 11000
ALLPIS = 207'b100001001100110111110011100100000010010111000001010010000010001001110000011111111110011101101110110100001111101000101111011010100101111101000010001101101111000010100110100110011011101000100000100110111100010;
XPCT = 108'b111100110101110100010000010010111100101101111101110101110000000010001110010000010011101010100111111010001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11200

pattern = 56; // 11200
ALLPIS = 207'b110000100110011011111001110010000001001011100000101001000001000100111000001111111111001110110111011010000111110100010111101101010010111110100001000110110111100001010011010011001101110100010000010011011110001;
XPCT = 108'b111010010110111010001000001011011110110011101111111111111001000111001110101100001001110100100001101101111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11400

pattern = 57; // 11400
ALLPIS = 207'b010001001101010011110001011001000100000010110011000110001000110010000110011010010110101001001001010011101111000001000001111100100110110100111011111110010100101010111111001000010010010100010101010001110000100;
XPCT = 108'b001001000001001010001010101001110000111010111001111110001111000010001111011100101010111111011000000111101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11600

pattern = 58; // 11600
ALLPIS = 207'b101000100110101001111000101100100010000001011001100011000100011001000011001101001011010100100100101001110111100000100000111110010011011010011101111111001010010101011111100100001001001010001010101000111000010;
XPCT = 108'b111100100100100101000101010100111000110011111110101111000000100011001010000000011100101011011110000001011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 11800

pattern = 59; // 11800
ALLPIS = 207'b010000001000101110101001110100000001110101100001110010100001100000100010100010100100000111111000000000101100011011110111000001111001101010111110011110011001011110000000100101110100110100100010101011000010110;
XPCT = 108'b000100101010011010010001010111000010101011111001111110010000100010111110011001101110100100111110110000001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12000

pattern = 60; // 12000
ALLPIS = 207'b101000010101001010000111010010000011010001110011011100010011110001010100010100011010001100001100000001001110111010010101100011001111100000100011110011111110010011000001011001010011110011010100000011100100110;
XPCT = 108'b110011000001111001101010000011100100111001101101111111111111011110001011100111000011111011111110100000011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12200

pattern = 61; // 12200
ALLPIS = 207'b111010011100100001011011101000100010101010111110100000100110011101110010100010101010101011001011000001100111000010111100011010111001000111001010011110010100000110110001111000001001100001010010111101111110010;
XPCT = 108'b110111000100110000101001011101111110010111111101011011111001000010000100000111110010111101100000101101000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12400

pattern = 62; // 12400
ALLPIS = 207'b111101001110010000101101110100010001010101011111010000010011001110111001010001010101010101100101100000110011100001011110001101011100100011100101001111001010000011011000111100000100110000101001011110111111001;
XPCT = 108'b110111100010011000010100101110111111100111111101111111010000110111011110110000100010101101011110001010101001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12600

pattern = 63; // 12600
ALLPIS = 207'b001111011011001010100010101001000101100000110110000110100101010011001100110110110001010010100001011000100000100011100000100010101110100010000111001101101011111110110110101010110101111000101000111100101101000;
XPCT = 108'b001101011010111100010100011100101101001101111001011010011111100000111111111101100110111000111001000000111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 12800

pattern = 64; // 12800
ALLPIS = 207'b110011111110011100000001011110010000101101101100010011001000110100010001101111001000010011010000010110100100010011001111001001010010000010011111101101000011100001101101001111011001101010101000100100001001100;
XPCT = 108'b110001110100110101010100010000001001011111111111011011000110110010011111011011111110100110011111101010111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13000

pattern = 65; // 13000
ALLPIS = 207'b011001111111001110000000101111001000010110110110001001100100011010001000110111100100001001101000001011010010001001100111100100101001000001001111110110100001110000110110100111101100110101010100010010000100110;
XPCT = 108'b001100111110011010101010001010000100100011111011111110001111011011101111001100010001110011000000101110100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13200

pattern = 66; // 13200
ALLPIS = 207'b001100101110111010010011111111100111100000011000100001110001001100000001011110111010001011000100000100110001110011011101110001100111110101011011000111100010000100011010011000011111110011101111011111000111110;
XPCT = 108'b001011000111111001110111101111000111101101111010101110000000100010000100011000100001101100011111000110101110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13400

pattern = 67; // 13400
ALLPIS = 207'b000110000110000000011010010111110000011011001111110101111011100111000101101010010101001010010010000011000000001110000000111011000000101111010001011111000011111110001100000111100110010000110010111001100110010;
XPCT = 108'b000000111011001000011001011101100110000011111010001010010110110000011011111001011101101101000111100010010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13600

pattern = 68; // 13600
ALLPIS = 207'b000011000011000000001101001011111000001101100111111010111101110011100010110101001010100101001001000001100000000111000000011101100000010111101000101111100001111111000110000011110011001000011001011100110011001;
XPCT = 108'b001000011001100100001100101100110011001111111001011010011111100011011111010111011101111111111110010011001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 13800

pattern = 69; // 13800
ALLPIS = 207'b100001110000111101010101001101111111101101110000011000011101111000110100011111101101011101010100100001101000110100001110001101000011011110001000101011000010000011100010001010010000001101001001111000011100001;
XPCT = 108'b111001010000000110100100111100011100101001111101110101111111111010011111100111000000110010000000011111111111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14000

pattern = 70; // 14000
ALLPIS = 207'b000111010001011111010001000011010110110110001100110001010010000100111010000100010001000110001110001010010111100110101011100011001110001010010011001110011111001111001001110111111100111101110000111011001000010;
XPCT = 108'b000110111110011110111000011111001000011001111010000000011111101100001111101111010001110001000001011101100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14200

pattern = 71; // 14200
ALLPIS = 207'b000011111001110010111011001001101000110000000101111101101010000011011000000111000000101100110111000100010011000100111011110010010100010000110101011011111101011011100101110000010111110111111101001011100001100;
XPCT = 108'b000110000011111011111110100111100001011011011011011010001111110000101111010100011011110000011000100110100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14400

pattern = 72; // 14400
ALLPIS = 207'b000001101101100100001110001100110111110011000001011011110110000000101001000110101000011001101011100011010001010101110011111010111001011101100110010001001100010001110011110011100010010010111011110011110101011;
XPCT = 108'b001110011001001001011101111011110101110011010011111110011111100100011111110100111110111000100000001111011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14600

pattern = 73; // 14600
ALLPIS = 207'b000000100111101111010100101110011000010010100011001000111000000001010001100110011100000011000101110000110000011101010111111110101111111011001111110100010100110100111000110010011000100000011000101111111111000;
XPCT = 108'b000110010100010000001100010111111111101101011000101110001111111011000101110110001010111110011111001011100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 14800

pattern = 74; // 14800
ALLPIS = 207'b100000010011110111101010010111001100001001010001100100011100000000101000110011001110000001100010111000011000001110101011111111010111111101100111111010001010011010011100011001001100010000001100010111111111100;
XPCT = 108'b110011000110001000000110001011111111100111111100101111011111011011111011011110010011111101011110000110100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15000

pattern = 75; // 15000
ALLPIS = 207'b000100010111010100111010000000111010110000111001010000110000010001010001010010000011111100000000010110001101111011100000111100110101011111001111001100101111000000010010111010011010010001010101100001011011001;
XPCT = 108'b001111010101001000101010110001011011101011111001111110001111011110101111010101000010111101011111000100111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15200

pattern = 76; // 15200
ALLPIS = 207'b000001000101110101001110100000001110101100001110010100001100000100010100010100100000111111000000000101100011011110111000001111001101010111110011110011001011110000000100101110100110100100010101011000010110110;
XPCT = 108'b000101111011010010001010101100010110100011111001111110001111011001001111011110100101111000000001011100000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15400

pattern = 77; // 15400
ALLPIS = 207'b000000100010111010100111010000000111010110000111001010000110000010001010001010010000011111100000000010110001101111011100000111100110101011111001111001100101111000000010010111010011010010001010101100001011011;
XPCT = 108'b001010110001101001000101010100001011101101111001111110000000100011010000010011111011101100000111000010010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15600

pattern = 78; // 15600
ALLPIS = 207'b111011100001101100011011101101101110110011001101011001000111010010001010111101010001111011111010111100011100011011001100011000100100100010110100000011001100111010000011000111100001111010000011100111111110000;
XPCT = 108'b111000111000111101000001110011111110010111111111011011111111100111001101011110011000111101011110011100001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 15800

pattern = 79; // 15800
ALLPIS = 207'b001011110100101111101011000100111000101110110100101110011111010111101011010100000101100000001011110010111100100101010010011101010001011101110000000101111011011010100110011100010100110010100110101100111110111;
XPCT = 108'b001011100010011001010011010100111110001111111001011010000000000110000100010000101010101101111001000100011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16000

pattern = 80; // 16000
ALLPIS = 207'b110111001000110110100101010000001010010100110110110000001011010001001101001001100111010100010010010010011100110001011101000000111010001001011011010000100011010010010001100010110000101000010001010100110001001;
XPCT = 108'b110100011000010100001000101000110001011111111101011011011111111100101111010101110011110001000000100010010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16200

pattern = 81; // 16200
ALLPIS = 207'b011101110010001101101001010100000010100101001101101100000010110100010011010010011001110101000100100100100111001100010111010000001110100010010110110100001000110100100100011000101100001010000100010101001100010;
XPCT = 108'b000011001110000101000010001001001100100111111001111110010000101110101110010011100011101011011110001100010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16400

pattern = 82; // 16400
ALLPIS = 207'b011000001001110000010101000010010011011100110010101110101101001101110100011011001001101011100100111000010001111011100100010000001101011100110000101010000000101101110110100000100010001010000010110010101001011;
XPCT = 108'b001100001001000101000001011010101001100011111001111110001111100100001111110101001110111011011110000011101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16600

pattern = 83; // 16600
ALLPIS = 207'b001001110001000101010101000000001101110001000010101100111010000010001101110001000010111001100010110010111011000101111011101111101000110000011111000100111101110010000011010101100100100001111001100110101010001;
XPCT = 108'b001010101010010000111100110010101010110101111001111110011111101000001111001100001101110011011001111011011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 16800

pattern = 84; // 16800
ALLPIS = 207'b011101111000000100101101101011100110011111111011111001001111110110011011110110110011110101110101010010111111110101110010001000100110010001011100011100000110010011100011010001110110001111001010101110110011010;
XPCT = 108'b001010001011000111100101010110110011111111000011111110010000111000111110000011001001100011011111111010011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17000

pattern = 85; // 17000
ALLPIS = 207'b101011001001111111001001010100110111010000100110000111001011011111111010000111111111110110101010000111101100000010110000100011111101010110101001011111111110101101001001101101001110100011011101101000100111001;
XPCT = 108'b110101100111010001101110110100100111010011111110000001011111111000111111110101111110111110111001011011100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17200

pattern = 86; // 17200
ALLPIS = 207'b011101111101011100000010000100101011100100111111100111101000000001010010100011001010110111110010011000010001000100100001011100100110000100101110101110111100111101110110011100011100111110010011111010001000000;
XPCT = 108'b001011100110011111001001111110001000101011111011111110011111101001001111111111100001110000011001101100110010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17400

pattern = 87; // 17400
ALLPIS = 207'b110001010101010101001111100000000111010011001010000001001011010010010001101010001010010000110110000100011011110100100000111000010011111111100110011101001001010101110010110001011001010101101110000000101110010;
XPCT = 108'b111110000100101010110111000000101110101011111111111111011111011100111111000100010111111110011111001001010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17600

pattern = 88; // 17600
ALLPIS = 207'b011101011111010111111000010001000111110110111110111011001001001101111111001001100011000100001011101100111110000010011001111011100111100001110100011111011001001110000001011101011001001110001111111111101001101;
XPCT = 108'b000011100100100111000111111111101001111111111011111110001111001001010011101110010001110011011000111100001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 17800

pattern = 89; // 17800
ALLPIS = 207'b101110101111101011111100001000100011111011011111011101100100100110111111100100110001100010000101110110011111000001001100111101110011110000111010001111101100100111000000101110101100100111000111111111110100110;
XPCT = 108'b110101111110010011100011111111110100000111111111010001000000110111101110110001000100100111011111011000001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18000

pattern = 90; // 18000
ALLPIS = 207'b010111010111110101111110000100010001111101101111101110110010010011011111110010011000110001000010111011001111100000100110011110111001111000011101000111110110010011100000010111010110010011100011111111111010011;
XPCT = 108'b000010110011001001110001111111111010001111111001011010010110000110101101010000011101100111111110111111011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18200

pattern = 91; // 18200
ALLPIS = 207'b001011101011111010111111000010001000111110110111110111011001001001101111111001001100011000100001011101100111110000010011001111011100111100001110100011111011001001110000001011101011001001110001111111111101001;
XPCT = 108'b000001011101100100111000111111111101000110101011011010011111010111101111000111110110111111111000011111010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18400

pattern = 92; // 18400
ALLPIS = 207'b110111100101001110101101101011101000110101011011101101001011100111101110001110011101011010110101111001010010101100000101010001001010001000111001000001011100100101010111000111100110000101000101110010001111100;
XPCT = 108'b111000111011000010100010111010001111010011111111011011101111110100111111010101110000110001011110000010110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18600

pattern = 93; // 18600
ALLPIS = 207'b011011110010100111010110110101110100011010101101110110100101110011110111000111001110101101011010111100101001010110000010101000100101000100011100100000101110010010101011100011110011000010100010111001000111110;
XPCT = 108'b001100011001100001010001011101000111011011111001011010000000000111001110010000011111101100000111110001101000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 18800

pattern = 94; // 18800
ALLPIS = 207'b111010011100011101000110110001010010111000001101010110011001011110010101101101111010001100011000100111000110000111000100000101011000101010110111010001001011101100000010110110011111100100010100101110101100011;
XPCT = 108'b111110110111110010001010010110101100001111111101011011110000000010101010011011001010100101000111001101111001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19000

pattern = 95; // 19000
ALLPIS = 207'b011001011000010111010101011001000100000000111010100111000100000001111110001001000110101010010100100110000101001101111011011100011100100011000100001010110000000110011110000100111001011111010001000000010001101;
XPCT = 108'b001000101100101111101000100000010001101011111011111110001111010011101101100111001010110101100000001100001011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19200

pattern = 96; // 19200
ALLPIS = 207'b100100101011101111111110001101001101001100000101000001010000111111001101001110011001011100100101000001111011010111010101101111011101100111010111111000001110110110011000100011011100010111110111010011010111001;
XPCT = 108'b110100010110001011111011101011010111101011110110101111111111100110111111010110111100110101011110001111100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19400

pattern = 97; // 19400
ALLPIS = 207'b111110101111110101010010001000111011100110011010111101011111101000011101011101111011001101111100101001001100011001110000001010111101010001001100111111011111001000110001001111010001000000111000000110111010010;
XPCT = 108'b110001110000100000011100000010111010011111011111011011100110111001110101100011100101101111111111001000111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19600

pattern = 98; // 19600
ALLPIS = 207'b010011011101010010110011011101001111000001101000110101110000000000000001111100110000101110100000111110110101000011010011010100100111011010010001001011100010011010101010000001110100110101000010101011011101100;
XPCT = 108'b001000001010011010100001010111011101001011111011011010001111101001001111111111010110110111011110000100100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 19800

pattern = 99; // 19800
ALLPIS = 207'b001000110001010011011110111000100110110001110101001010000101110100011001001010101010010110110010000100000110010000000001011111000110000010010001000011100101110011001001110000010110101110001101001110011110101;
XPCT = 108'b000110000011010111000110100110011110111111111000101110001111001000100101000101111010110010011111000100011111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20000

pattern = 100; // 20000
ALLPIS = 207'b110011111101100111000010110111111011101101100001001000001001011101100010101011001000010001101100111011010001100100000101111110101001001001110001100000101110011100110011111111101101010010000011010101000000110;
XPCT = 108'b111111111110101001000001101001000000010111111101011011000110110011101111111011011001101001011111101010110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20200

pattern = 101; // 20200
ALLPIS = 207'b011101101101001011101110100011001011000111000001111111100100111000011011010010010111101111010111011011110011011010100010000111010000001101010010101100101011100001001101111100001110101000110010100011101111110;
XPCT = 108'b000111100111010100011001010011101111110011111011111110001111111010001111100111110000111010000110101101100010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20400

pattern = 102; // 20400
ALLPIS = 207'b111001010011101011011010111010001101010110111011010010111001111011100011100111010110101101011110010100101011000001010100010010100010001110010000010111001001010101110001111001100001010001011100100011111000011;
XPCT = 108'b110111001000101000101110010011111000110011111101111111111111011000001111111111011011111010011001000111110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20600

pattern = 103; // 20600
ALLPIS = 207'b001110000101000010100110101111001110011101100000110011111101010100101010111011001100001111001100110101100011000101000001000111101010101001011111001001110110110011101011010110010011101011011010101111011101011;
XPCT = 108'b001010110001110101101101010111011101011101111010001010000000000111111110100001111001101010111110110111011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 20800

pattern = 104; // 20800
ALLPIS = 207'b011100001100010110001001010000111100000111001100010111001011011001000011000001100010011011000010001010001101011011101000110101100100110010000001000001100011011000111011101000111100111011101101001111001111011;
XPCT = 108'b001101001110011101110110100111001111111111111011111110000000101101101110001011100100101000011110011011110001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21000

pattern = 105; // 21000
ALLPIS = 207'b010001101011101110001011010010001001100110110011011011101010010100101011010100110101110101100010010101100010101011000101011011001000001001010011000000101110000010110101100110000100001010011111000000101011010;
XPCT = 108'b000100110010000101001111100000101011110011111011111110011111001101001111100100100001111111000001100111010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21200

pattern = 106; // 21200
ALLPIS = 207'b010010110010010000001011110010100100111110101100101000100010000111110001010001100000001110001010010010011001010111001110000000100011000111100111100000111101010100010110000101101010000110000011100011010010010;
XPCT = 108'b001000101101000011000001110011010010000010111001011010010110010100001111111001001111100111011110110110000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21400

pattern = 107; // 21400
ALLPIS = 207'b101110100101010110011110010100100101011110110110110110100101001100000101110000010010001101110010000110011011110100011000010111000111111111000110011001011101010010000110100110101101000111001111110110010110111;
XPCT = 108'b111100111110100011100111111010010110000111111101011011110110111111001111011010001110100111011111100111111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21600

pattern = 108; // 21600
ALLPIS = 207'b101010001010111010010001100001101001110000000111100110001000101110111001001011010100110100101101110000011111011111110101100100010001011100110100001101101101001110110111000010110001001001000100110110001001101;
XPCT = 108'b111000011000100100100010011010001001011101111101010001001111000100100101100101011111111011100001010000011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 21800

pattern = 109; // 21800
ALLPIS = 207'b110110010001011001000001100110111101000100001110010111010011100000101111001010110011011101001011001001011110000100001100011101011100110010110101011001001110000111110000011000001111111101110011000100010110000;
XPCT = 108'b110011000111111110111001100000010110000111110111011011101111011001011111100111110001111111111110001101000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22000

pattern = 110; // 22000
ALLPIS = 207'b110111101010011110100011111110100100101010011011100101001110110001001001110000111111010100110011110110010011001010011110110100010111111100110000011110111011001100011000111100011000000101011111101010100111000;
XPCT = 108'b110111100100000010101111110110100111001010111111011011010000110101001110000011010100101011011111001001110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22200

pattern = 111; // 22200
ALLPIS = 207'b010101010000100001001001101000110001101001110001101110101110110010000110100101010000011110110010001011011101100111110100001000010001101111101110001001010011000001010101011001101010011010010110100101001000111;
XPCT = 108'b000011001101001101001011010001001000110111111001111110001001011101101010011110110001111110000000111011111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22400

pattern = 112; // 22400
ALLPIS = 207'b100100001010011000010101110111001100001010101101011101010000001001100011010000010011010110010101011000010001010000101001011000000011010000010011010111001001010101110111111111000100001001110000100001011110111;
XPCT = 108'b111111110010000100111000010001011110110001111111111111010110110101001111001010000000101011000110101001010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22600

pattern = 113; // 22600
ALLPIS = 207'b001111010011111111000100111011001110000110100101000000000111100010110111111110110111101000101110011111011010010000000110001011011100000110110001101100111100010010101101100111111110111111101111001100000001101;
XPCT = 108'b000100111111011111110111100100000001011101111000000000001111010111011111100111111110110000011001011111001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 22800

pattern = 114; // 22800
ALLPIS = 207'b011001000101100100000110011011110100010000111001011101001110000010111100101011001101110100101100100101111000010000110001110101110011001011010101100100111000011111000001100000111111110111001100010001011000001;
XPCT = 108'b000100001111111011100110001001011000111011111011111110011111001010011011011111101001110000111111001010000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23000

pattern = 115; // 23000
ALLPIS = 207'b110001011001011100101111111111111101100110100100010001011100001111111110101011110101010010011000101000100000110110110001010011101111001110001110101111000000101110011010011110000111010000011100000000010110010;
XPCT = 108'b111011110011101000001110000000010110100011111111111111010000111100011110101001111010101100111110111010011010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23200

pattern = 116; // 23200
ALLPIS = 207'b010110111100000000000000101010101011001110101000101101000000011011010101101100001101100100011011011101011011101011011001000100111000111100001011101111000111100000000101011001110010001010001000011111110000111;
XPCT = 108'b000011001001000101000100001111110000011111111011011010001111001100111111000101110001111011000000110000110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23400

pattern = 117; // 23400
ALLPIS = 207'b100011110010001000100001011011001111011111010000100001010101110111100000100101110101110010001101001011101011010111100100001101100010110011110110000010000011100011110000100011111001010111010000110011111110100;
XPCT = 108'b110100011100101011101000011011111110001001110111011011001001000100101110101110111100111100000000011000011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23600

pattern = 118; // 23600
ALLPIS = 207'b001111001011100100000000000010111111001101010101001011001100000001000001001000000110111110100010101000111011011101000111010100111101101101000100110000100101111100111001100110100100011011000000010011110100101;
XPCT = 108'b000100111010001101100000001011110100010001111010001010001111110011111111101101001100111010111000000000010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 23800

pattern = 119; // 23800
ALLPIS = 207'b101101000110100011001100110011100001110100000101000110101001100110001000110001000101111000001000001010100100100101000101100011000011010110001001101010100011010010000110000001101111111001010101010001111010100;
XPCT = 108'b111000001111111100101010101001111010100011111101111111100000100000101110010001101111101000111111100000000010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24000

pattern = 120; // 24000
ALLPIS = 207'b111011010001101000110011001100111000011101000001010001101010011001100010001100010001011110000010000010101001001001010001011000110000110101100010011010101000110100100001100000011011111110010101010100011110101;
XPCT = 108'b110100000101111111001010101000011110011111111111011011101111101010001111010101000010110001011110001001011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24200

pattern = 121; // 24200
ALLPIS = 207'b011110110011110010101101101001110000110111110000010011101100110010100001110101011011001000101101000011011100011110110010100000010011010100111011010111011001010100001110110000010100011011011111110111110000101;
XPCT = 108'b001110000010001101101111111011110000001111111011011010001111000000111111011100001000111010111000010100010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24400

pattern = 122; // 24400
ALLPIS = 207'b000000110111010000001100100101011000100111101011010100110001100110001101101011111001110011100001001100011110000111101011101110000100011000101000111100101011111000011011000100110000111111011011101001100100001;
XPCT = 108'b001000101000011111101101110101100100111011110000101110001111111101101111000111111111110000011111100100011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24600

pattern = 123; // 24600
ALLPIS = 207'b110110001100010001100011001110001101100000000100011101111100000111010111000011101101100010000111010001100110111110000000100101101101010110100000101111011110110101011011101101101101111000100110010001111011111;
XPCT = 108'b111101101110111100010011001001111011010011101111011011000000100001011110100011110100100111011110101010010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 24800

pattern = 124; // 24800
ALLPIS = 207'b011100110110011100011000111111001000110000000111000000100100101111111000011101010010011001000101010110110100010010010101101001101101000110101111001110100010110100011011111000111000100011000001110110100001001;
XPCT = 108'b001111001100010001100000111010100001111111111001111110000000010110011110101000100010101111011110110011110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25000

pattern = 125; // 25000
ALLPIS = 207'b101001101011011010100101000111101010011000000110101110001000111011101111110010001101100100100100010101011101000100011111001111101101001110101000111110011100110100111011110010010010001110110010000101001100010;
XPCT = 108'b111110010001000111011001000001001100111100111100101111011001000000101100100110000100111100000111100000011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25200

pattern = 126; // 25200
ALLPIS = 207'b110011101010000111000111011101011101000010001011101100011001110111110011110011110101001100000111001001110000101101001111110100000101111110110001111110100101001100001000100100010111111110111101101100001000100;
XPCT = 108'b110100100011111111011110110100001000001111111101011011101001110111011110101101101010111111000001101011001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25400

pattern = 127; // 25400
ALLPIS = 207'b011111001010110111110111010001111010001011001011101100111111011011110000111000111011110110001110100101111000001010010010101001111111110010111001011010110010101001110110000001111101100011101010100000110110000;
XPCT = 108'b001000001110110001110101010000110110001011111001011010010000001101011100111001111111101110111111110111000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25600

pattern = 128; // 25600
ALLPIS = 207'b011001100110001101101010111001111101011011100110011110011111000111100111011101010001010111100100101010110110001000110110000100100100011010000110010111010000110100101110110010110101100001010100110100101100000;
XPCT = 108'b001110011010110000101010011000101100101111111001111110011111100101101101001101110011110011000000010011001000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 25800

pattern = 129; // 25800
ALLPIS = 207'b001011110101101111111010101111110100011100011000110101001110101001100101001101010001101000111000101000001010000101111011000111001000010000100011001000000001000000000011011000001011000110011101111101111111010;
XPCT = 108'b001011000101100011001110111101111111010111111011011010011001000101010110000101000011111100011001001110000110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26000

pattern = 130; // 26000
ALLPIS = 207'b010001101010010001111100110010001100000111111010110110000101011110111011011111000111001000010011110110111101010001111000000000101010011111111101011110100101010001101010010001101110010111011000100001001000100;
XPCT = 108'b001010001111001011101100010001001000100011011001111110001001101100001110101100001011110010100001100010010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26200

pattern = 131; // 26200
ALLPIS = 207'b001111111111001101111011101100100101101001000111111101110111010010111101011100000001110010000101010111011010000010111001111010010110101000100100110001010110001110110111100011111110111110000011000101001000010;
XPCT = 108'b001100011111011111000001100001001000011111111011010000011111110101010011001110101100110000100001110000111010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26400

pattern = 132; // 26400
ALLPIS = 207'b100111000010001101111101100000001011100001011011000010110111000000110011111000011100111011111000001011101000011100011000011111101100000011001011101111100001110011010000001011111101001011110011111100010000010;
XPCT = 108'b110001011110100101111001111100010000001111111101010001110000111101111100011000010011101101111000110111011110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26600

pattern = 133; // 26600
ALLPIS = 207'b010001100000011100010000110100011110000010101011001111100011001011001011010100010100001101111010110110000000011000011110110011101100011101010001000110000100011011100110100100011000000000110011101100111000100;
XPCT = 108'b001100100100000000011001110100111000101111111011111110001111100010101111101100100010110001000001001001000000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 26800

pattern = 134; // 26800
ALLPIS = 207'b011001011001010000001010011100111010100101110101100100110000010011000100000000101000010011010110000101111000101001010010111111100101001100000101100111110000101100010001010001011100000101011011111011101000010;
XPCT = 108'b000010000110000010101101111111101000111011111001111110011111010100111111101101001011111010111001111010011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27000

pattern = 135; // 27000
ALLPIS = 207'b010011001110110000111011100111111101010000110001101110100011110011111100100010101110100110101110101100001100111111100100010001010110010010000001001110000101000100011111000100110000011000010001000101100011010;
XPCT = 108'b001000101000001100001000100001100011011111111001011010010000000100101100011011010111100100111110111100011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27200

pattern = 136; // 27200
ALLPIS = 207'b010000110111111111110110100000100110100010011100100010110111010110110000000000001010000001010100010010011010100001111001110111001101000100110001001110000110100110010110111100000001000111011010011000000110000;
XPCT = 108'b001111100000100011101101001100000110100011111001111110011111011111010101010100000010110111011111000000101100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27400

pattern = 137; // 27400
ALLPIS = 207'b111001110011011001111011101100110111000001010001011100110111001011010111011000100110111101011000001000100000100011011110111010011001011110001111100010101111011000010001110001000111010000000110111001011101011;
XPCT = 108'b110110000011101000000011011101011101110011111101111111111111111111111111101110000010111111011111000001010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27600

pattern = 138; // 27600
ALLPIS = 207'b100111001100110110111111010010001011010011000100001011011111001011110101111100000000101111001010100111100001100101100110111000010111110001110111110010001000111010010011001011000000011001110000001011100000100;
XPCT = 108'b111001010000001100111000000111100000010011111111010001100000011100111110111000001100101010011111011111000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 27800

pattern = 139; // 27800
ALLPIS = 207'b000010000011101001011011001111001000010100101001111000101100000100000010111010100101010011010111010111100110101100101110110110100101110111000101011100000101001000011010101101011010011011010000001011011001101;
XPCT = 108'b001101100101001101101000000111011001001011111000001010001111111000111111010100110110111001011110000000010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28000

pattern = 140; // 28000
ALLPIS = 207'b101001110111011001110101111010010101110100100001110011010011011100000000111010011010101111101111001101001000101110010000100001001010110010111100101111101110000101011000001100100110110011010010001110111010110;
XPCT = 108'b110001101011011001101001000110111010100101111110101111101111001101111111011101000001110110011000010110100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28200

pattern = 141; // 28200
ALLPIS = 207'b111010010101110100010010001011010000011010111100110011110000010100011010110010010000010000110011001111000001011101011001011010111001111010010100100100011111100110110101111100001001101100100010110001001000101;
XPCT = 108'b110111100100110110010001011001001000010010110111011011011111100101111111100100110000110010011110000110111011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28400

pattern = 142; // 28400
ALLPIS = 207'b100001011110001110001101100110101101111011001010110001110110101011000111001111110100001110001101001101000111101010110100110100101000011001000110011101110111010111010110000111110010101111100000000100111101110;
XPCT = 108'b111000111001010111110000000000111101101111011111111111100000011011011110100011110010100001100110000111011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28600

pattern = 143; // 28600
ALLPIS = 207'b110101001110011101011100011011101101100011011111001100011000011011011110101111010110010010001100011111101101101111011111111111101110110001010110011000000100111011111010100111100111101101010001001010001000001;
XPCT = 108'b111100111011110110101000100110001000100011011101111111011111100000011111101110000100111111000000111100010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 28800

pattern = 144; // 28800
ALLPIS = 207'b011010100111001110101110001101110110110001101111100110001100001101101111010111101011001001000110001111110110110111101111111111110111011000101011001100000010011101111101010011110011110110101000100101000100000;
XPCT = 108'b000010011001111011010100010001000100011111101001011010011111011010011111101100101011110100111111001110100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29000

pattern = 145; // 29000
ALLPIS = 207'b000101111011000010011011101100011000111111110001100000100110110111100110110000101001101111111001111000001011110101110101001001010011100100011111000100111010100110001100110111011011001000100011011100101110111;
XPCT = 108'b000110110101100100010001101100101110101111111000101110000110010111111111101010111100101101111111111010001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29200

pattern = 146; // 29200
ALLPIS = 207'b011011101100110100001111011000000101011110110100111100100000110100111011110111111111101110101110101011111100101010101110101000101111001000010100100100111101101001101001110110101000010111010011110111101100101;
XPCT = 108'b000110111100001011101001111011101100010111111001011010000110011101111111111011011011100101011111100111011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29400

pattern = 147; // 29400
ALLPIS = 207'b010000111011101011111000110001110000100110101110011110111001100111110000111101111010011111110010101000001101110110101000111011101001011111000101000001010000010110000000111101101011100110011101011011011001111;
XPCT = 108'b000111101101110011001110101111011001100011111001111110011111000101011111111110110010110101011000000000010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29600

pattern = 148; // 29600
ALLPIS = 207'b011100010101000010100010100010001010100111111111010101100101110000101001001010111010000111000011101111011010110111110000101011111111010000010000000001000001101010001111001110010011101110010000011011011110101;
XPCT = 108'b001001110001110111001000001111011110111011111011111110001111000000001111000110010101110010111000111101000111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 29800

pattern = 149; // 29800
ALLPIS = 207'b100001100001111101110011010101110001011000100000100101101110011001110100000101000001010000010000110111100111100011011011011010010111000001100010100100000011100100111011100110010111110001110001110001100000010;
XPCT = 108'b111100110011111000111000111001100000111001111110100101011001000000001110111100100010110000000001110100111000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30000

pattern = 150; // 30000
ALLPIS = 207'b110001001000101100101110110101110110001001011001110001111000010110010001100100110001100111111100101101001101111001101010110001010000011111100010001111101100100100010111111000100100011011111001101110010001100;
XPCT = 108'b111111001010001101111100110110010001110111111111111111000110110110111111000011111110101100011110101000010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30200

pattern = 151; // 30200
ALLPIS = 207'b111101101100100111010010111101011110011100000001100101101100100010001101110100100011000001011001010100100010101101101011001110101010101111110101100011000111001001010100111000001000101001011100110111010110010;
XPCT = 108'b110111000100010100101110011011010110100111111111111111010000101011111110111000010000101011011110111111100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30400

pattern = 152; // 30400
ALLPIS = 207'b001011101110011001001100011011010110000111101111110010010110101011001010010000011111111010001011010111000110011001011101000101011000010001010011010011100011010100111111100001000101101010100011110101100111101;
XPCT = 108'b001100000010110101010001111001100111010111111000001010001111001111101111100101000011111100000001100111011001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30600

pattern = 153; // 30600
ALLPIS = 207'b001000010110000010011110100001110000000100110100001001001111101000010001101100100011000010110111000111001110011010010010010100010110100001100110011001011100100011100010000011001001111100100111011010001010111;
XPCT = 108'b001000010100111110010011101110001010100011111011111110000000100101001110110000011101100000111000011011010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 30800

pattern = 154; // 30800
ALLPIS = 207'b101000010001111101001001011110001001001001101100111101001101011110111101101110011011011100100000101110010000111010111000000110000100011111000101000010101101111010011110001000101011000111100000111110111010111;
XPCT = 108'b111001001101100011110000011110111010100111011110100101101111000100101111011100100101110111011110010111110011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31000

pattern = 155; // 31000
ALLPIS = 207'b110110111000010011100111101111010110001101111110101000111101011011001111111001110001010100100110110101100000101101010101111010010100010100001011011101100000100111111100011000111010000011110000000010010001110;
XPCT = 108'b110011001101000001111000000010010001001011111101011011011001001100111110110110010011111111100001100111100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31200

pattern = 156; // 31200
ALLPIS = 207'b111001000100111000011010010000111011000000011100011011101000010101000000001111001001010001011001010101101101011010100100111101100010010001111000100100110010001110100101001111100100110110100101101110100111100;
XPCT = 108'b110001111010011011010010110110100111110111111111111111000110010100101001010001111100100001011111111001110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31400

pattern = 157; // 31400
ALLPIS = 207'b010101111000100111100010001100100110000101010100110111010010001000010011111111011010100101110000000011000001011101011010010011100101111001000101110001110101110100101101011110111101001010110100001100011110001;
XPCT = 108'b000011111110100101011010000100011110111111011011111110010000100001100110100011100110101000111111000111101111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31600

pattern = 158; // 31600
ALLPIS = 207'b110101110010000000000100010111110100101110011111000000010100011011110011011000110100111101101010000010011000010001010100111101111000011010101010110110000110010101101011111100110001000010100001001110011001001;
XPCT = 108'b111111101000100001010000100110011001111111111101111111110110001101111111010011001100100010011111101000100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 31800

pattern = 159; // 31800
ALLPIS = 207'b100100111010000101010001001001111001000101101010011110010101101111101001111010110001011010111001001001001110010010001111001100100101011001110000000010111100100011011001000001111100110011111011101010110111000;
XPCT = 108'b110000001110011001111101110110110111111001111100101111101111011110001111100110101111111100000001010111001010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32000

pattern = 160; // 32000
ALLPIS = 207'b100110101100111000000000000010010101100110100000111111001010011110101011100001000000100100001101110111111011000001011111111111000100001100001011000000001100000000010110010100010111100010010011100111110100110;
XPCT = 108'b111010100011110001001001110011110100001101111111011011010000101101111110010000001001101110011110000000000100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32200

pattern = 161; // 32200
ALLPIS = 207'b111110000001111010010111000010101000111011100001101100110000100000110111010101011010110101000101001111111111110100011110111000000011010001011111100101111101000010010101111000111110001001000100111111001011100;
XPCT = 108'b110111001111000100100010011111001011011110000101011011001111100010110101000110110010111011011000101001111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32400

pattern = 162; // 32400
ALLPIS = 207'b010111110101100011100010101000000010111110101000100110101010001011101110001100100111110011101101000100010000000001111000010100110000110101101110001111001011100101010011111000111101000011111001110000001000110;
XPCT = 108'b001111001110100001111100111000001000011011111001011010001111111011111111001111001001110001011001111011100000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32600

pattern = 163; // 32600
ALLPIS = 207'b100011000001110000011101100011001101000101001001010100110011011110101010000101110010101101001110111100110100000011111000110010000000000110110001101100010101010001011010101010111011010110001011001010011111111;
XPCT = 108'b111101011101101011000101100110011111001011111100001011101111110100011111010101000001111100000110011011100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 32800

pattern = 164; // 32800
ALLPIS = 207'b110001100000111000001110110001100110100010100100101010011001101111010101000010111001010110100111011110011010000001111100011001000000000011011000110110001010101000101101010101011101101011000101100101001111111;
XPCT = 108'b110010100110110101100010110001001111111111111101111111000110000001000111010011011000100101011110100010001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33000

pattern = 165; // 33000
ALLPIS = 207'b111011101011100110110001000110010001001010011100010110000100101111101010111011000101011110101110011010001000101001011100010100010001001011100101010010101100111110010011110000101100011001111100011001110110110;
XPCT = 108'b111110001110001100111110001101110110010011111101011011101111111110101111010100101000110110111110011111001110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33200

pattern = 166; // 33200
ALLPIS = 207'b011100011111000011001010100001100101010101111110100010101100001011001000000000111100100000110000010000101101111111000011001001010001011011110000111101111111111110001101000000100111010111001100110100111111110;
XPCT = 108'b000000001011101011100110011000111111110111111001111110011111111001101111100101011111110101011000111101100110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33400

pattern = 167; // 33400
ALLPIS = 207'b100011100001100001011111000110001011001110100010011101110111100111000000001111101001111011010010100001110011001010001001000010001100101111100001111010110101111111101100101001111101000111001110001110110001100;
XPCT = 108'b110101001110100011100111000110110001001111111110001011101111001101101111110111010011110101111111100111010110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33600

pattern = 168; // 33600
ALLPIS = 207'b111011101110110100101011011010010010011100011111111101001011110000110100110100011111110010111110110110111001000010000110100101001110010011001100011000110000100000010101110000001010111110101101001000101000101;
XPCT = 108'b110110000101011111010110100100101000010010111111011011001001001111111110001110100100110010000000100000000011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 33800

pattern = 169; // 33800
ALLPIS = 207'b110100000001000000000001101111011010011110010100110100000110010000111110110000010100011110011100001011101010100001001111100110110110011110110101100110001000100010011000100001111101100100001011100101010100100;
XPCT = 108'b110100001110110010000101110001010100101111111101111111101111110000000101010100101110110110011111000010101010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34000

pattern = 170; // 34000
ALLPIS = 207'b101001100010011010000011001010111101110100111101111100101110110011100110000101101100001011110001011101100101111010010010001101001000011111101001010000101011111011011011000011100011011010011001110111110000010;
XPCT = 108'b111000011001101101001100111011110000110101111100101111110000010000011110011000001101100000011000001010010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34200

pattern = 171; // 34200
ALLPIS = 207'b011111001100000101100110000000100001000011100001100111101001100101010001011001010111001010111011000101110000101001000110011100101101011101111110100111110000101100101110010110000111010000000011001101100010101;
XPCT = 108'b001010110011101000000001100101100010000111111011011010000000110011111110111010011001101101111110000011010011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34400

pattern = 172; // 34400
ALLPIS = 207'b100100010111000001011000110010100000100101100010110011000101011001000011001010001100001100111111010111101010000011111010111011100111011001110001101001110000001111110011011011110011010100000010110110101101100;
XPCT = 108'b111011011001101010000001011010101101111111111111111111101111101001000101000111010001110100111110000100010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34600

pattern = 173; // 34600
ALLPIS = 207'b001110100000111011000001111000111001101011100111111011000100100010001100010111100010011000011110101001011111100100100011001101110111100011100100100100000110011001000111000000000110001000010101111110101100101;
XPCT = 108'b001000000011000100001010111110101100010101111011011010010000001001001110100011101101101011011110101110100001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 34800

pattern = 174; // 34800
ALLPIS = 207'b001001001100111001110100000001001110111110000011101101000101110101100110100110101011011110011000110010110001111100101110011010101010000111111100000010101101011010110001100010101011010111101101100010000111001;
XPCT = 108'b000100011101101011110110110010000111110001111011111110011111110011101111100111011011111111000000001001010111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35000

pattern = 175; // 35000
ALLPIS = 207'b011101101100011000100011101001001111110010000010010110100011110001010110100100100010111110010010011111101101001010100101110000110110100101011011110011000001110101101100000110000110000000100111010010101001100;
XPCT = 108'b000000110011000000010011101010101001100011111001111110000110110010111111011011001111101111011111110010110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35200

pattern = 176; // 35200
ALLPIS = 207'b111011000010000000011010000000010110110010110110000010000101110101100110011100010110110010001010010101001111100110000000011011101000110010010100101110011110000001000101100011101011010101110111000110101001100;
XPCT = 108'b110100011101101010111011100010101001010111011101011011001001011001001110010110010111110110100001000100111100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35400

pattern = 177; // 35400
ALLPIS = 207'b001111001011100000100000010010001000100110101101111100011110101100011001010100101111100111001101100111100011110000011110111011010000011011010011101000100000111011010100110001000000001101100001011001111000101;
XPCT = 108'b000110000000000110110000101101111000000001111001011010001111101010011111010101111010110100111001001110011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35600

pattern = 178; // 35600
ALLPIS = 207'b101101011000101010111100100110111100100010011111011010111111001111110010010011000110111101101011010000000111000010001110000000111010001010111101111010000111011110000000000010001110000000111101010101111111100;
XPCT = 108'b110000010111000000011110101001111111100111111101110101100000111100101110110011101111101111011111100011110000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 35800

pattern = 179; // 35800
ALLPIS = 207'b011001000110010011110011111011100001011010010011101011010110101010011011110001111101010100010100101010101110101000111101110100101011110101011110101111101110010011111111000101000001110110010100001100111000001;
XPCT = 108'b001000100000111011001010000100111000110111111011111110011001100010001110011101010010111100000000011100111101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36000

pattern = 180; // 36000
ALLPIS = 207'b010010100000111101011111001011011011101011001101001001110111000000011011111011010111001111100110011001001010111011100100100101001111011000101110100001011110000000000011001110000111001001110110011100110110110;
XPCT = 108'b001001110011100100111011001100110110010111111011011010000000100101101110100000000101101011000111100010110110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36200

pattern = 181; // 36200
ALLPIS = 207'b011111100101000010110110010000101111101011111011100011001010111010111101000000011011111011111000110111100111011101111110101001110111111010010101111101110000110010001110100111111100010000100000000101111110010;
XPCT = 108'b001100111110001000010000000001111110001111111011011010010110000000110011011011111100101101111111110111100100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36400

pattern = 182; // 36400
ALLPIS = 207'b111011011010100100100011100110001000000000110100101000010000100111101001100110000011011011100010111111111111100001110101001100101100000011001011011010010110001010010100111111011001110110101101011010101110111;
XPCT = 108'b110111110100111011010110101110101110001011111101011011100000110111011110110010011110101100000000101011001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36600

pattern = 183; // 36600
ALLPIS = 207'b010110001001001000001001110010000001011000111010010111010110111111101101001111111000010100010001011101101000110101101100111101100000010101111001000011011111001111000011101101000000000010110011011011100010101;
XPCT = 108'b001101100000000001011001101111100010010011110011011010001111011001001111100111100100111111111110111110010101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 36800

pattern = 184; // 36800
ALLPIS = 207'b101100000010000010100011011100101110101101111111100010111101110000000101110100000100101000001010100000000100011111010001101100111110001101000011101001001011101001110111110110101011110111110011110101000101101;
XPCT = 108'b111110111101111011111001111001000101110101111101111111110000010000010100000001101010100100111111101011001101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37000

pattern = 185; // 37000
ALLPIS = 207'b001000100011001100010001011110101010000000010111111000111000011111101010001100011101010110100011001100000001101011011110110000001101110010110100110010101110010101110010011000101001101000010000000111001000001;
XPCT = 108'b001011001100110100001000000011001000100101011001111110011111000101111111011100110011111010011111100010010001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37200

pattern = 186; // 37200
ALLPIS = 207'b011101011110100001101111111010000110111010101001010010000010101100110111101110000001111011110101101000100000100001100101001111010010100100100011101111001101010110110110000000000100000010000100010110100101101;
XPCT = 108'b001000000010000001000010001010100101100111111001111110000000111011001010110011111111101111011111001010000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37400

pattern = 187; // 37400
ALLPIS = 207'b011110001010101010110011100011011001010000011010000000101001011010000100100111111000011100010111010111101000001010111001000010000010110111111011110110110001001001100111111011010000100011111111111100110101001;
XPCT = 108'b001111010000010001111111111100110101011111111001011010010000000100101110100000000010101111111111111111000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37600

pattern = 188; // 37600
ALLPIS = 207'b111100011011011011001011111000000010010000011001100101110001011100110101000010111101011000101101111001010110011101111011011110000101001000101100001110111010100001011100101000111010101111100011111000000001111;
XPCT = 108'b110101001101010111110001111100000001101011110111111111111111000111011011010111010100110010011001100100110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 37800

pattern = 189; // 37800
ALLPIS = 207'b000000001111111011001010110110101111100000011110001101011100001011110110100010111100001110111111000011001100101101100010111011111001101001111100101011000110000001011000101100000011111100111010000001011000000;
XPCT = 108'b000101100001111110011101000001011000100011111010100100001111101010011111100111010100111111011110011001010010;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38000

pattern = 190; // 38000
ALLPIS = 207'b110110010110000100111000001001000010100110100100011011011000100011011101010011000101001100100011000010010110011111000000101110011000100111110111001010000000001010101110110000000011111001101001010001100000101;
XPCT = 108'b111110000001111100110100101001100000000011111111011011111111010010011111010100111000111000100001100111001111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38200

pattern = 191; // 38200
ALLPIS = 207'b100100110010001110000011000011010111010000010100000111101111011100001100101100000010111100000001101010001010001100111011111010010011011000001000010000001101100011001110101000010100010000111100111100000111010;
XPCT = 108'b111101000010001000011110011100000111101101110110101111111001111011111110110110100100111101100001011111111110;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38400

pattern = 192; // 38400
ALLPIS = 207'b101000111100101001101000101001011111011000100110110101001110111000111000101001011111100011101101110101001101010110111000100010001001100001000011101110001010100100001110101110000011011111100000110011000101010;
XPCT = 108'b111101110001101111110000011011000101100011111110100101010000010111000000110000000100100001000111011000010000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38600

pattern = 193; // 38600
ALLPIS = 207'b010101010001100000011110101011111101001011001100100111011011000010111101100000000100001111111000110110010111001000000011100111001111001110101100101110110010011100000001101100101011111011000110011101110100111;
XPCT = 108'b000101101101111101100011001101110100110111111011111110001111010000001111000101111110111000000110000000011101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 38800

pattern = 194; // 38800
ALLPIS = 207'b011101000100011110100111101100010000001011001101000000011010110011011000111001100111000100000001101010110001010110111011100111000110100000100010010110110010100100101100000010101101000011001111010110011000101;
XPCT = 108'b000000011110100001100111101010011000100111111001111110000000100011101110111011001111101111011111100011100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39000

pattern = 195; // 39000
ALLPIS = 207'b000100100110001001010110000011100001111101000000010100000000110111111111111010011000100001000000010010011010010000111101010000111101111110001111001101011101100101100000001001011110110010100100111100110111001;
XPCT = 108'b000001000111011001010010011100110111101101111001110100011111101000101111110101110111111100000001110110011011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39200

pattern = 196; // 39200
ALLPIS = 207'b010110000100111100000100010010001011000110001000100111000001001000110011100111101001010011010011110110000100010011011111100010101011101010100100110100111000100100010011110010111011001001000101101000010011101;
XPCT = 108'b001110011101100100100010110100010011011011111011011010001001000000101110100111001000111010000000100101000001;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39400

pattern = 197; // 39400
ALLPIS = 207'b111110010100110011101011111011000110010010111111011001111110100110101111001011011111111100011000000000100110000111000000011000100000011000000011101100101110101111100101011001111100100001001110011111110101000;
XPCT = 108'b110011001110010000100111001111110101011111111111011011110000010111001110001000110001101111011110011111110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39600

pattern = 198; // 39600
ALLPIS = 207'b001000101010010101011101000011110101011100101000101000000001111010100011000011101111010000101001111111000011100100010001001100000001001000100010000100101100001011110110110001110111000001001001010011110000001;
XPCT = 108'b001110001011100000100100101011110000101011110001111110001111000010001111111110111010111110000000110110000101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 39800

pattern = 199; // 39800
ALLPIS = 207'b001100101010100101001011010010001000000111010101001100010010110101000001000001001011101111111011001100111110100100010001011011000001000011100010011011100110001101101101011000001111110010110101001010110001110;
XPCT = 108'b000011000111111001011010100110110001110011111000101110010000101010101110100000100011101100111110100110011100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40000

pattern = 200; // 40000
ALLPIS = 207'b000010101111011110100000000111101101110000110101010100101010101010111110101011010000000101111111001101101111011000101110111010100111111010001001011010001101101111011111100100101100000110100100010100011011000;
XPCT = 108'b001100101110000011010010001000011011010101111000000000011111101100011111101110101110110111111110101001010100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40200

pattern = 201; // 40200
ALLPIS = 207'b110011011110011111110110000011010001111100101110100011111100001111000011111100001010101111010110010011000101110110011110011110001101010001111001001110111111100011001011001001110000011011010001001110100000100;
XPCT = 108'b111001001000001101101000100110100000011111111111011011100000000111001110001010101100101010011111001010011000;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40400

pattern = 202; // 40400
ALLPIS = 207'b111001000111001000100111100001101111110110011010100010001011110001111110110010101101010011101001010000100000100011010101101011010000010011110000001100010101010111001111001011101001101011001001101010101011001;
XPCT = 108'b111001011100110101100100110110101011110011111101111111011111001011111111111100110110110101111110110001100011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40600

pattern = 203; // 40600
ALLPIS = 207'b010101100101001111111110110011101000101110111110010100100000110100001011111011110110101011100011101001110111110101111010110011101111011110011100101001101000111011000111010111111000111001010111101001011110010;
XPCT = 108'b001010111100011100101011110101011110111011101001111110011111000011001111110101000100111000000001111101001100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 40800

pattern = 204; // 40800
ALLPIS = 207'b100000000010010000111011010001101100110001111000101000000001001011000000011110010101011010011001110110101001001110101110101011100100101010000110010011001000110110101111010101000110110101001111001000000101011;
XPCT = 108'b111010100011011010100111100100000101110011110100101111100000001111111110101000011011100100111110100111100111;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41000

pattern = 205; // 41000
ALLPIS = 207'b010100010011111011110110100011011100001100010000010000000001011101010101100111110000110010000101011101000010011101011110111101001011100001101001000011111011010011111011000010111110100000111001110001010100011;
XPCT = 108'b001000011111010000011100111001010100111011110001111110001001101101101110000101001111111110000110100011110101;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41200

pattern = 206; // 41200
ALLPIS = 207'b100101010011111001110000010010001000011011100011100101100100000100000000011110001010001011110001000000100010000110100111110010000111111011011110100011000001101100010001000101010100010111010100101011100101111;
XPCT = 108'b110000100010001011101010010111100101111001111111111111101111001000101111110101111010111110111001100111101011;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41400

pattern = 207; // 41400
ALLPIS = 207'b000100101101111100010110001101000100101010000101001011100010000111011001010001000100000010100001000011011000000110110101101010111100110000000001000001011111010011100100001101011011100001001101111011110110100;
XPCT = 108'b000001100101110000100110111111110110101001111011111110001111000110011111110100000101111110111111001011110100;
MASK = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#0 ->capture;
#200; // 41600

      $display("// %t : Simulation of %0d patterns completed with %0d errors\n", $time, pattern+1, nofails);
      if (verbose >=2) $finish(2);
      /* else */ $finish(0);
   end
endmodule
