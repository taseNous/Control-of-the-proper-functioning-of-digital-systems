`ifndef __FIFO_TB__
`define __FIFO_TB__
//-----------------------------------------------------------------------------
`include "fifo.v"
`include "fifo_property.sv"
`include "fifo_test.sv"
`include "fifo_if.sv"
//-----------------------------------------------------------------------------
`define DUV   duv
//-----------------------------------------------------------------------------
module fifo_tb;
//-----------------------------------------------------------------------------
bit clk, rstn;
//-----------------------------------------------------------------------------
localparam  fifo_depth = 8;
localparam  fifo_width = 8;
//-----------------------------------------------------------------------------
clkrstn_if clkrstn();
fifo_if #(.dw(fifo_width)) fwrite_if (.clk(clk),.rstn(rstn));
fifo_if #(.dw(fifo_width)) fread_if  (.clk(clk),.rstn(rstn));
//-----------------------------------------------------------------------------
/**
 * Clock
 */
always #5 clk=!clk;
//-----------------------------------------------------------------------------
initial begin : reset
    rstn = 1'b0;
    repeat(2) begin @(posedge clk); end
    #2 rstn = 1'b1;
end
//-----------------------------------------------------------------------------
assign clkrstn.clk  = clk;
assign clkrstn.rstn = rstn;
//-----------------------------------------------------------------------------
fifo_test oop_tb (
//-----------------------------------------------------------------------------
    .clkrstn    ( clkrstn   ),
    .fifo_read  ( fread_if  ),
    .fifo_write ( fwrite_if )
);
//-----------------------------------------------------------------------------
/**
 * Device-Under-Verification
 */
//-----------------------------------------------------------------------------
fifo #(
//-----------------------------------------------------------------------------
    .fifo_depth     ( fifo_depth    ),
    .fifo_width     ( fifo_width    )
//-----------------------------------------------------------------------------
  ) duv (
//-----------------------------------------------------------------------------
    .clk            ( clk            ),
    .rstn           ( rstn           ),
    //---------------------------------
    .fifo_data_out  ( fread_if.data  ),
    .fifo_empty     ( fread_if.req   ),
    .fifo_read      ( fread_if.ack   ),
    //---------------------------------
    .fifo_data_in   ( fwrite_if.data ),
    .fifo_full      ( fwrite_if.ack  ),
    .fifo_write     ( fwrite_if.req  )
    //---------------------------------
);
//-----------------------------------------------------------------------------
/**
 * Bind checker
 */
//-----------------------------------------------------------------------------
bind `DUV fifo_property#(
//-----------------------------------------------------------------------------
    .fifo_depth(fifo_depth),
    .fifo_width(fifo_width)
//-----------------------------------------------------------------------------
  ) duv_bind (
//-----------------------------------------------------------------------------
    .clk            ( clk           ),
    .rstn           ( rstn          ),
    .fifo_data_out  ( fifo_data_out ),
    .fifo_full      ( fifo_full     ),
    .fifo_empty     ( fifo_empty    ),
    .fifo_write     ( fifo_write    ),
    .fifo_read      ( fifo_read     ),
    .fifo_data_in   ( fifo_data_in  )
);
//-----------------------------------------------------------------------------
endmodule
//-----------------------------------------------------------------------------
`endif