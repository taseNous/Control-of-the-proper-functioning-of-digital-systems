`ifndef __GEN_CLS__
`define __GEN_CLS__
//------------------------------------------------------------------------------
`include "dat_cls.svh"
//------------------------------------------------------------------------------
class gen_cls /*#(int data_width = 8)*/;
//------------------------------------------------------------------------------

    // Transaction
    //-------------------------------------
    dat_cls rngdat;
    //-------------------------------------
    integer cnt;

    // Mailbox
    //-------------------------------------
    mailbox mbox;

    // Constructor
    //-------------------------------------
    function new(mailbox mbox, integer cnt);
        this.mbox = mbox;
        this.cnt  = cnt;
    endfunction : new
    //-------------------------------------

    // Main Task
    //-------------------------------------
    task main();
    //-------------------------------------
        repeat(cnt) begin
            rngdat = new();
            if(!rngdat.randomize()) begin
                $fatal(1,"[fatal]: unable to generate transtaction");
            end
            rngdat.show("gen");
            mbox.put(rngdat);
        end
    //-------------------------------------
    endtask
    //-------------------------------------

//------------------------------------------------------------------------------
endclass: gen_cls
//------------------------------------------------------------------------------
`endif